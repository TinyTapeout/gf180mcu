magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< psubdiff >>
rect 0 69943 400 69968
rect 0 69871 130 69943
rect 0 69825 25 69871
rect 71 69825 130 69871
rect 0 69803 130 69825
rect 270 69871 400 69943
rect 270 69825 329 69871
rect 375 69825 400 69871
rect 270 69803 400 69825
rect 0 69778 400 69803
rect 0 69708 93 69778
rect 0 13356 25 69708
rect 71 13356 93 69708
rect 307 69708 400 69778
rect 0 13287 93 13356
rect 307 13356 329 69708
rect 375 13356 400 69708
rect 307 13287 400 13356
rect 0 13262 400 13287
rect 0 13231 130 13262
rect 0 13185 25 13231
rect 71 13185 130 13231
rect 0 13122 130 13185
rect 270 13231 400 13262
rect 270 13185 329 13231
rect 375 13185 400 13231
rect 270 13122 400 13185
rect 0 13097 400 13122
<< psubdiffcont >>
rect 25 69825 71 69871
rect 130 69803 270 69943
rect 329 69825 375 69871
rect 25 13356 71 69708
rect 329 13356 375 69708
rect 25 13185 71 13231
rect 130 13122 270 13262
rect 329 13185 375 13231
<< polysilicon >>
rect 155 69687 239 69706
rect 155 69641 174 69687
rect 220 69641 239 69687
rect 155 69527 239 69641
rect 155 69481 174 69527
rect 220 69481 239 69527
rect 155 69367 239 69481
rect 155 69321 174 69367
rect 220 69321 239 69367
rect 155 69207 239 69321
rect 155 69161 174 69207
rect 220 69161 239 69207
rect 155 69047 239 69161
rect 155 69001 174 69047
rect 220 69001 239 69047
rect 155 68887 239 69001
rect 155 68841 174 68887
rect 220 68841 239 68887
rect 155 68727 239 68841
rect 155 68681 174 68727
rect 220 68681 239 68727
rect 155 68567 239 68681
rect 155 68521 174 68567
rect 220 68521 239 68567
rect 155 68407 239 68521
rect 155 68361 174 68407
rect 220 68361 239 68407
rect 155 68247 239 68361
rect 155 68201 174 68247
rect 220 68201 239 68247
rect 155 68087 239 68201
rect 155 68041 174 68087
rect 220 68041 239 68087
rect 155 67927 239 68041
rect 155 67881 174 67927
rect 220 67881 239 67927
rect 155 67767 239 67881
rect 155 67721 174 67767
rect 220 67721 239 67767
rect 155 67607 239 67721
rect 155 67561 174 67607
rect 220 67561 239 67607
rect 155 67447 239 67561
rect 155 67401 174 67447
rect 220 67401 239 67447
rect 155 67287 239 67401
rect 155 67241 174 67287
rect 220 67241 239 67287
rect 155 67127 239 67241
rect 155 67081 174 67127
rect 220 67081 239 67127
rect 155 66967 239 67081
rect 155 66921 174 66967
rect 220 66921 239 66967
rect 155 66807 239 66921
rect 155 66761 174 66807
rect 220 66761 239 66807
rect 155 66647 239 66761
rect 155 66601 174 66647
rect 220 66601 239 66647
rect 155 66487 239 66601
rect 155 66441 174 66487
rect 220 66441 239 66487
rect 155 66327 239 66441
rect 155 66281 174 66327
rect 220 66281 239 66327
rect 155 66167 239 66281
rect 155 66121 174 66167
rect 220 66121 239 66167
rect 155 66007 239 66121
rect 155 65961 174 66007
rect 220 65961 239 66007
rect 155 65847 239 65961
rect 155 65801 174 65847
rect 220 65801 239 65847
rect 155 65687 239 65801
rect 155 65641 174 65687
rect 220 65641 239 65687
rect 155 65527 239 65641
rect 155 65481 174 65527
rect 220 65481 239 65527
rect 155 65367 239 65481
rect 155 65321 174 65367
rect 220 65321 239 65367
rect 155 65207 239 65321
rect 155 65161 174 65207
rect 220 65161 239 65207
rect 155 65047 239 65161
rect 155 65001 174 65047
rect 220 65001 239 65047
rect 155 64887 239 65001
rect 155 64841 174 64887
rect 220 64841 239 64887
rect 155 64727 239 64841
rect 155 64681 174 64727
rect 220 64681 239 64727
rect 155 64567 239 64681
rect 155 64521 174 64567
rect 220 64521 239 64567
rect 155 64407 239 64521
rect 155 64361 174 64407
rect 220 64361 239 64407
rect 155 64247 239 64361
rect 155 64201 174 64247
rect 220 64201 239 64247
rect 155 64087 239 64201
rect 155 64041 174 64087
rect 220 64041 239 64087
rect 155 63927 239 64041
rect 155 63881 174 63927
rect 220 63881 239 63927
rect 155 63767 239 63881
rect 155 63721 174 63767
rect 220 63721 239 63767
rect 155 63607 239 63721
rect 155 63561 174 63607
rect 220 63561 239 63607
rect 155 63447 239 63561
rect 155 63401 174 63447
rect 220 63401 239 63447
rect 155 63287 239 63401
rect 155 63241 174 63287
rect 220 63241 239 63287
rect 155 63127 239 63241
rect 155 63081 174 63127
rect 220 63081 239 63127
rect 155 62967 239 63081
rect 155 62921 174 62967
rect 220 62921 239 62967
rect 155 62807 239 62921
rect 155 62761 174 62807
rect 220 62761 239 62807
rect 155 62647 239 62761
rect 155 62601 174 62647
rect 220 62601 239 62647
rect 155 62487 239 62601
rect 155 62441 174 62487
rect 220 62441 239 62487
rect 155 62327 239 62441
rect 155 62281 174 62327
rect 220 62281 239 62327
rect 155 62167 239 62281
rect 155 62121 174 62167
rect 220 62121 239 62167
rect 155 62007 239 62121
rect 155 61961 174 62007
rect 220 61961 239 62007
rect 155 61847 239 61961
rect 155 61801 174 61847
rect 220 61801 239 61847
rect 155 61687 239 61801
rect 155 61641 174 61687
rect 220 61641 239 61687
rect 155 61527 239 61641
rect 155 61481 174 61527
rect 220 61481 239 61527
rect 155 61367 239 61481
rect 155 61321 174 61367
rect 220 61321 239 61367
rect 155 61207 239 61321
rect 155 61161 174 61207
rect 220 61161 239 61207
rect 155 61047 239 61161
rect 155 61001 174 61047
rect 220 61001 239 61047
rect 155 60887 239 61001
rect 155 60841 174 60887
rect 220 60841 239 60887
rect 155 60727 239 60841
rect 155 60681 174 60727
rect 220 60681 239 60727
rect 155 60567 239 60681
rect 155 60521 174 60567
rect 220 60521 239 60567
rect 155 60407 239 60521
rect 155 60361 174 60407
rect 220 60361 239 60407
rect 155 60247 239 60361
rect 155 60201 174 60247
rect 220 60201 239 60247
rect 155 60087 239 60201
rect 155 60041 174 60087
rect 220 60041 239 60087
rect 155 59927 239 60041
rect 155 59881 174 59927
rect 220 59881 239 59927
rect 155 59767 239 59881
rect 155 59721 174 59767
rect 220 59721 239 59767
rect 155 59607 239 59721
rect 155 59561 174 59607
rect 220 59561 239 59607
rect 155 59447 239 59561
rect 155 59401 174 59447
rect 220 59401 239 59447
rect 155 59287 239 59401
rect 155 59241 174 59287
rect 220 59241 239 59287
rect 155 59127 239 59241
rect 155 59081 174 59127
rect 220 59081 239 59127
rect 155 58967 239 59081
rect 155 58921 174 58967
rect 220 58921 239 58967
rect 155 58807 239 58921
rect 155 58761 174 58807
rect 220 58761 239 58807
rect 155 58647 239 58761
rect 155 58601 174 58647
rect 220 58601 239 58647
rect 155 58487 239 58601
rect 155 58441 174 58487
rect 220 58441 239 58487
rect 155 58327 239 58441
rect 155 58281 174 58327
rect 220 58281 239 58327
rect 155 58167 239 58281
rect 155 58121 174 58167
rect 220 58121 239 58167
rect 155 58007 239 58121
rect 155 57961 174 58007
rect 220 57961 239 58007
rect 155 57847 239 57961
rect 155 57801 174 57847
rect 220 57801 239 57847
rect 155 57687 239 57801
rect 155 57641 174 57687
rect 220 57641 239 57687
rect 155 57527 239 57641
rect 155 57481 174 57527
rect 220 57481 239 57527
rect 155 57367 239 57481
rect 155 57321 174 57367
rect 220 57321 239 57367
rect 155 57207 239 57321
rect 155 57161 174 57207
rect 220 57161 239 57207
rect 155 57047 239 57161
rect 155 57001 174 57047
rect 220 57001 239 57047
rect 155 56887 239 57001
rect 155 56841 174 56887
rect 220 56841 239 56887
rect 155 56727 239 56841
rect 155 56681 174 56727
rect 220 56681 239 56727
rect 155 56567 239 56681
rect 155 56521 174 56567
rect 220 56521 239 56567
rect 155 56407 239 56521
rect 155 56361 174 56407
rect 220 56361 239 56407
rect 155 56247 239 56361
rect 155 56201 174 56247
rect 220 56201 239 56247
rect 155 56087 239 56201
rect 155 56041 174 56087
rect 220 56041 239 56087
rect 155 55927 239 56041
rect 155 55881 174 55927
rect 220 55881 239 55927
rect 155 55767 239 55881
rect 155 55721 174 55767
rect 220 55721 239 55767
rect 155 55607 239 55721
rect 155 55561 174 55607
rect 220 55561 239 55607
rect 155 55447 239 55561
rect 155 55401 174 55447
rect 220 55401 239 55447
rect 155 55287 239 55401
rect 155 55241 174 55287
rect 220 55241 239 55287
rect 155 55127 239 55241
rect 155 55081 174 55127
rect 220 55081 239 55127
rect 155 54967 239 55081
rect 155 54921 174 54967
rect 220 54921 239 54967
rect 155 54807 239 54921
rect 155 54761 174 54807
rect 220 54761 239 54807
rect 155 54647 239 54761
rect 155 54601 174 54647
rect 220 54601 239 54647
rect 155 54487 239 54601
rect 155 54441 174 54487
rect 220 54441 239 54487
rect 155 54327 239 54441
rect 155 54281 174 54327
rect 220 54281 239 54327
rect 155 54167 239 54281
rect 155 54121 174 54167
rect 220 54121 239 54167
rect 155 54007 239 54121
rect 155 53961 174 54007
rect 220 53961 239 54007
rect 155 53847 239 53961
rect 155 53801 174 53847
rect 220 53801 239 53847
rect 155 53687 239 53801
rect 155 53641 174 53687
rect 220 53641 239 53687
rect 155 53527 239 53641
rect 155 53481 174 53527
rect 220 53481 239 53527
rect 155 53367 239 53481
rect 155 53321 174 53367
rect 220 53321 239 53367
rect 155 53207 239 53321
rect 155 53161 174 53207
rect 220 53161 239 53207
rect 155 53047 239 53161
rect 155 53001 174 53047
rect 220 53001 239 53047
rect 155 52887 239 53001
rect 155 52841 174 52887
rect 220 52841 239 52887
rect 155 52727 239 52841
rect 155 52681 174 52727
rect 220 52681 239 52727
rect 155 52567 239 52681
rect 155 52521 174 52567
rect 220 52521 239 52567
rect 155 52407 239 52521
rect 155 52361 174 52407
rect 220 52361 239 52407
rect 155 52247 239 52361
rect 155 52201 174 52247
rect 220 52201 239 52247
rect 155 52087 239 52201
rect 155 52041 174 52087
rect 220 52041 239 52087
rect 155 51927 239 52041
rect 155 51881 174 51927
rect 220 51881 239 51927
rect 155 51767 239 51881
rect 155 51721 174 51767
rect 220 51721 239 51767
rect 155 51607 239 51721
rect 155 51561 174 51607
rect 220 51561 239 51607
rect 155 51447 239 51561
rect 155 51401 174 51447
rect 220 51401 239 51447
rect 155 51287 239 51401
rect 155 51241 174 51287
rect 220 51241 239 51287
rect 155 51127 239 51241
rect 155 51081 174 51127
rect 220 51081 239 51127
rect 155 50967 239 51081
rect 155 50921 174 50967
rect 220 50921 239 50967
rect 155 50807 239 50921
rect 155 50761 174 50807
rect 220 50761 239 50807
rect 155 50647 239 50761
rect 155 50601 174 50647
rect 220 50601 239 50647
rect 155 50487 239 50601
rect 155 50441 174 50487
rect 220 50441 239 50487
rect 155 50327 239 50441
rect 155 50281 174 50327
rect 220 50281 239 50327
rect 155 50167 239 50281
rect 155 50121 174 50167
rect 220 50121 239 50167
rect 155 50007 239 50121
rect 155 49961 174 50007
rect 220 49961 239 50007
rect 155 49847 239 49961
rect 155 49801 174 49847
rect 220 49801 239 49847
rect 155 49687 239 49801
rect 155 49641 174 49687
rect 220 49641 239 49687
rect 155 49527 239 49641
rect 155 49481 174 49527
rect 220 49481 239 49527
rect 155 49367 239 49481
rect 155 49321 174 49367
rect 220 49321 239 49367
rect 155 49207 239 49321
rect 155 49161 174 49207
rect 220 49161 239 49207
rect 155 49047 239 49161
rect 155 49001 174 49047
rect 220 49001 239 49047
rect 155 48887 239 49001
rect 155 48841 174 48887
rect 220 48841 239 48887
rect 155 48727 239 48841
rect 155 48681 174 48727
rect 220 48681 239 48727
rect 155 48567 239 48681
rect 155 48521 174 48567
rect 220 48521 239 48567
rect 155 48407 239 48521
rect 155 48361 174 48407
rect 220 48361 239 48407
rect 155 48247 239 48361
rect 155 48201 174 48247
rect 220 48201 239 48247
rect 155 48087 239 48201
rect 155 48041 174 48087
rect 220 48041 239 48087
rect 155 47927 239 48041
rect 155 47881 174 47927
rect 220 47881 239 47927
rect 155 47767 239 47881
rect 155 47721 174 47767
rect 220 47721 239 47767
rect 155 47607 239 47721
rect 155 47561 174 47607
rect 220 47561 239 47607
rect 155 47447 239 47561
rect 155 47401 174 47447
rect 220 47401 239 47447
rect 155 47287 239 47401
rect 155 47241 174 47287
rect 220 47241 239 47287
rect 155 47127 239 47241
rect 155 47081 174 47127
rect 220 47081 239 47127
rect 155 46967 239 47081
rect 155 46921 174 46967
rect 220 46921 239 46967
rect 155 46807 239 46921
rect 155 46761 174 46807
rect 220 46761 239 46807
rect 155 46647 239 46761
rect 155 46601 174 46647
rect 220 46601 239 46647
rect 155 46487 239 46601
rect 155 46441 174 46487
rect 220 46441 239 46487
rect 155 46327 239 46441
rect 155 46281 174 46327
rect 220 46281 239 46327
rect 155 46167 239 46281
rect 155 46121 174 46167
rect 220 46121 239 46167
rect 155 46007 239 46121
rect 155 45961 174 46007
rect 220 45961 239 46007
rect 155 45847 239 45961
rect 155 45801 174 45847
rect 220 45801 239 45847
rect 155 45687 239 45801
rect 155 45641 174 45687
rect 220 45641 239 45687
rect 155 45527 239 45641
rect 155 45481 174 45527
rect 220 45481 239 45527
rect 155 45367 239 45481
rect 155 45321 174 45367
rect 220 45321 239 45367
rect 155 45207 239 45321
rect 155 45161 174 45207
rect 220 45161 239 45207
rect 155 45047 239 45161
rect 155 45001 174 45047
rect 220 45001 239 45047
rect 155 44887 239 45001
rect 155 44841 174 44887
rect 220 44841 239 44887
rect 155 44727 239 44841
rect 155 44681 174 44727
rect 220 44681 239 44727
rect 155 44567 239 44681
rect 155 44521 174 44567
rect 220 44521 239 44567
rect 155 44407 239 44521
rect 155 44361 174 44407
rect 220 44361 239 44407
rect 155 44247 239 44361
rect 155 44201 174 44247
rect 220 44201 239 44247
rect 155 44087 239 44201
rect 155 44041 174 44087
rect 220 44041 239 44087
rect 155 43927 239 44041
rect 155 43881 174 43927
rect 220 43881 239 43927
rect 155 43767 239 43881
rect 155 43721 174 43767
rect 220 43721 239 43767
rect 155 43607 239 43721
rect 155 43561 174 43607
rect 220 43561 239 43607
rect 155 43447 239 43561
rect 155 43401 174 43447
rect 220 43401 239 43447
rect 155 43287 239 43401
rect 155 43241 174 43287
rect 220 43241 239 43287
rect 155 43127 239 43241
rect 155 43081 174 43127
rect 220 43081 239 43127
rect 155 42967 239 43081
rect 155 42921 174 42967
rect 220 42921 239 42967
rect 155 42807 239 42921
rect 155 42761 174 42807
rect 220 42761 239 42807
rect 155 42647 239 42761
rect 155 42601 174 42647
rect 220 42601 239 42647
rect 155 42487 239 42601
rect 155 42441 174 42487
rect 220 42441 239 42487
rect 155 42327 239 42441
rect 155 42281 174 42327
rect 220 42281 239 42327
rect 155 42167 239 42281
rect 155 42121 174 42167
rect 220 42121 239 42167
rect 155 42007 239 42121
rect 155 41961 174 42007
rect 220 41961 239 42007
rect 155 41847 239 41961
rect 155 41801 174 41847
rect 220 41801 239 41847
rect 155 41687 239 41801
rect 155 41641 174 41687
rect 220 41641 239 41687
rect 155 41527 239 41641
rect 155 41481 174 41527
rect 220 41481 239 41527
rect 155 41367 239 41481
rect 155 41321 174 41367
rect 220 41321 239 41367
rect 155 41207 239 41321
rect 155 41161 174 41207
rect 220 41161 239 41207
rect 155 41047 239 41161
rect 155 41001 174 41047
rect 220 41001 239 41047
rect 155 40887 239 41001
rect 155 40841 174 40887
rect 220 40841 239 40887
rect 155 40727 239 40841
rect 155 40681 174 40727
rect 220 40681 239 40727
rect 155 40567 239 40681
rect 155 40521 174 40567
rect 220 40521 239 40567
rect 155 40407 239 40521
rect 155 40361 174 40407
rect 220 40361 239 40407
rect 155 40247 239 40361
rect 155 40201 174 40247
rect 220 40201 239 40247
rect 155 40087 239 40201
rect 155 40041 174 40087
rect 220 40041 239 40087
rect 155 39927 239 40041
rect 155 39881 174 39927
rect 220 39881 239 39927
rect 155 39767 239 39881
rect 155 39721 174 39767
rect 220 39721 239 39767
rect 155 39607 239 39721
rect 155 39561 174 39607
rect 220 39561 239 39607
rect 155 39447 239 39561
rect 155 39401 174 39447
rect 220 39401 239 39447
rect 155 39287 239 39401
rect 155 39241 174 39287
rect 220 39241 239 39287
rect 155 39127 239 39241
rect 155 39081 174 39127
rect 220 39081 239 39127
rect 155 38967 239 39081
rect 155 38921 174 38967
rect 220 38921 239 38967
rect 155 38807 239 38921
rect 155 38761 174 38807
rect 220 38761 239 38807
rect 155 38647 239 38761
rect 155 38601 174 38647
rect 220 38601 239 38647
rect 155 38487 239 38601
rect 155 38441 174 38487
rect 220 38441 239 38487
rect 155 38327 239 38441
rect 155 38281 174 38327
rect 220 38281 239 38327
rect 155 38167 239 38281
rect 155 38121 174 38167
rect 220 38121 239 38167
rect 155 38007 239 38121
rect 155 37961 174 38007
rect 220 37961 239 38007
rect 155 37847 239 37961
rect 155 37801 174 37847
rect 220 37801 239 37847
rect 155 37687 239 37801
rect 155 37641 174 37687
rect 220 37641 239 37687
rect 155 37527 239 37641
rect 155 37481 174 37527
rect 220 37481 239 37527
rect 155 37367 239 37481
rect 155 37321 174 37367
rect 220 37321 239 37367
rect 155 37207 239 37321
rect 155 37161 174 37207
rect 220 37161 239 37207
rect 155 37047 239 37161
rect 155 37001 174 37047
rect 220 37001 239 37047
rect 155 36887 239 37001
rect 155 36841 174 36887
rect 220 36841 239 36887
rect 155 36727 239 36841
rect 155 36681 174 36727
rect 220 36681 239 36727
rect 155 36567 239 36681
rect 155 36521 174 36567
rect 220 36521 239 36567
rect 155 36407 239 36521
rect 155 36361 174 36407
rect 220 36361 239 36407
rect 155 36247 239 36361
rect 155 36201 174 36247
rect 220 36201 239 36247
rect 155 36087 239 36201
rect 155 36041 174 36087
rect 220 36041 239 36087
rect 155 35927 239 36041
rect 155 35881 174 35927
rect 220 35881 239 35927
rect 155 35767 239 35881
rect 155 35721 174 35767
rect 220 35721 239 35767
rect 155 35607 239 35721
rect 155 35561 174 35607
rect 220 35561 239 35607
rect 155 35447 239 35561
rect 155 35401 174 35447
rect 220 35401 239 35447
rect 155 35287 239 35401
rect 155 35241 174 35287
rect 220 35241 239 35287
rect 155 35127 239 35241
rect 155 35081 174 35127
rect 220 35081 239 35127
rect 155 34967 239 35081
rect 155 34921 174 34967
rect 220 34921 239 34967
rect 155 34807 239 34921
rect 155 34761 174 34807
rect 220 34761 239 34807
rect 155 34647 239 34761
rect 155 34601 174 34647
rect 220 34601 239 34647
rect 155 34487 239 34601
rect 155 34441 174 34487
rect 220 34441 239 34487
rect 155 34327 239 34441
rect 155 34281 174 34327
rect 220 34281 239 34327
rect 155 34167 239 34281
rect 155 34121 174 34167
rect 220 34121 239 34167
rect 155 34007 239 34121
rect 155 33961 174 34007
rect 220 33961 239 34007
rect 155 33847 239 33961
rect 155 33801 174 33847
rect 220 33801 239 33847
rect 155 33687 239 33801
rect 155 33641 174 33687
rect 220 33641 239 33687
rect 155 33527 239 33641
rect 155 33481 174 33527
rect 220 33481 239 33527
rect 155 33367 239 33481
rect 155 33321 174 33367
rect 220 33321 239 33367
rect 155 33207 239 33321
rect 155 33161 174 33207
rect 220 33161 239 33207
rect 155 33047 239 33161
rect 155 33001 174 33047
rect 220 33001 239 33047
rect 155 32887 239 33001
rect 155 32841 174 32887
rect 220 32841 239 32887
rect 155 32727 239 32841
rect 155 32681 174 32727
rect 220 32681 239 32727
rect 155 32567 239 32681
rect 155 32521 174 32567
rect 220 32521 239 32567
rect 155 32407 239 32521
rect 155 32361 174 32407
rect 220 32361 239 32407
rect 155 32247 239 32361
rect 155 32201 174 32247
rect 220 32201 239 32247
rect 155 32087 239 32201
rect 155 32041 174 32087
rect 220 32041 239 32087
rect 155 31927 239 32041
rect 155 31881 174 31927
rect 220 31881 239 31927
rect 155 31767 239 31881
rect 155 31721 174 31767
rect 220 31721 239 31767
rect 155 31607 239 31721
rect 155 31561 174 31607
rect 220 31561 239 31607
rect 155 31447 239 31561
rect 155 31401 174 31447
rect 220 31401 239 31447
rect 155 31287 239 31401
rect 155 31241 174 31287
rect 220 31241 239 31287
rect 155 31127 239 31241
rect 155 31081 174 31127
rect 220 31081 239 31127
rect 155 30967 239 31081
rect 155 30921 174 30967
rect 220 30921 239 30967
rect 155 30807 239 30921
rect 155 30761 174 30807
rect 220 30761 239 30807
rect 155 30647 239 30761
rect 155 30601 174 30647
rect 220 30601 239 30647
rect 155 30487 239 30601
rect 155 30441 174 30487
rect 220 30441 239 30487
rect 155 30327 239 30441
rect 155 30281 174 30327
rect 220 30281 239 30327
rect 155 30167 239 30281
rect 155 30121 174 30167
rect 220 30121 239 30167
rect 155 30007 239 30121
rect 155 29961 174 30007
rect 220 29961 239 30007
rect 155 29847 239 29961
rect 155 29801 174 29847
rect 220 29801 239 29847
rect 155 29687 239 29801
rect 155 29641 174 29687
rect 220 29641 239 29687
rect 155 29527 239 29641
rect 155 29481 174 29527
rect 220 29481 239 29527
rect 155 29367 239 29481
rect 155 29321 174 29367
rect 220 29321 239 29367
rect 155 29207 239 29321
rect 155 29161 174 29207
rect 220 29161 239 29207
rect 155 29047 239 29161
rect 155 29001 174 29047
rect 220 29001 239 29047
rect 155 28887 239 29001
rect 155 28841 174 28887
rect 220 28841 239 28887
rect 155 28727 239 28841
rect 155 28681 174 28727
rect 220 28681 239 28727
rect 155 28567 239 28681
rect 155 28521 174 28567
rect 220 28521 239 28567
rect 155 28407 239 28521
rect 155 28361 174 28407
rect 220 28361 239 28407
rect 155 28247 239 28361
rect 155 28201 174 28247
rect 220 28201 239 28247
rect 155 28087 239 28201
rect 155 28041 174 28087
rect 220 28041 239 28087
rect 155 27927 239 28041
rect 155 27881 174 27927
rect 220 27881 239 27927
rect 155 27767 239 27881
rect 155 27721 174 27767
rect 220 27721 239 27767
rect 155 27607 239 27721
rect 155 27561 174 27607
rect 220 27561 239 27607
rect 155 27447 239 27561
rect 155 27401 174 27447
rect 220 27401 239 27447
rect 155 27287 239 27401
rect 155 27241 174 27287
rect 220 27241 239 27287
rect 155 27127 239 27241
rect 155 27081 174 27127
rect 220 27081 239 27127
rect 155 26967 239 27081
rect 155 26921 174 26967
rect 220 26921 239 26967
rect 155 26807 239 26921
rect 155 26761 174 26807
rect 220 26761 239 26807
rect 155 26647 239 26761
rect 155 26601 174 26647
rect 220 26601 239 26647
rect 155 26487 239 26601
rect 155 26441 174 26487
rect 220 26441 239 26487
rect 155 26327 239 26441
rect 155 26281 174 26327
rect 220 26281 239 26327
rect 155 26167 239 26281
rect 155 26121 174 26167
rect 220 26121 239 26167
rect 155 26007 239 26121
rect 155 25961 174 26007
rect 220 25961 239 26007
rect 155 25847 239 25961
rect 155 25801 174 25847
rect 220 25801 239 25847
rect 155 25687 239 25801
rect 155 25641 174 25687
rect 220 25641 239 25687
rect 155 25527 239 25641
rect 155 25481 174 25527
rect 220 25481 239 25527
rect 155 25367 239 25481
rect 155 25321 174 25367
rect 220 25321 239 25367
rect 155 25207 239 25321
rect 155 25161 174 25207
rect 220 25161 239 25207
rect 155 25047 239 25161
rect 155 25001 174 25047
rect 220 25001 239 25047
rect 155 24887 239 25001
rect 155 24841 174 24887
rect 220 24841 239 24887
rect 155 24727 239 24841
rect 155 24681 174 24727
rect 220 24681 239 24727
rect 155 24567 239 24681
rect 155 24521 174 24567
rect 220 24521 239 24567
rect 155 24407 239 24521
rect 155 24361 174 24407
rect 220 24361 239 24407
rect 155 24247 239 24361
rect 155 24201 174 24247
rect 220 24201 239 24247
rect 155 24087 239 24201
rect 155 24041 174 24087
rect 220 24041 239 24087
rect 155 23927 239 24041
rect 155 23881 174 23927
rect 220 23881 239 23927
rect 155 23767 239 23881
rect 155 23721 174 23767
rect 220 23721 239 23767
rect 155 23607 239 23721
rect 155 23561 174 23607
rect 220 23561 239 23607
rect 155 23447 239 23561
rect 155 23401 174 23447
rect 220 23401 239 23447
rect 155 23287 239 23401
rect 155 23241 174 23287
rect 220 23241 239 23287
rect 155 23127 239 23241
rect 155 23081 174 23127
rect 220 23081 239 23127
rect 155 22967 239 23081
rect 155 22921 174 22967
rect 220 22921 239 22967
rect 155 22807 239 22921
rect 155 22761 174 22807
rect 220 22761 239 22807
rect 155 22647 239 22761
rect 155 22601 174 22647
rect 220 22601 239 22647
rect 155 22487 239 22601
rect 155 22441 174 22487
rect 220 22441 239 22487
rect 155 22327 239 22441
rect 155 22281 174 22327
rect 220 22281 239 22327
rect 155 22167 239 22281
rect 155 22121 174 22167
rect 220 22121 239 22167
rect 155 22007 239 22121
rect 155 21961 174 22007
rect 220 21961 239 22007
rect 155 21847 239 21961
rect 155 21801 174 21847
rect 220 21801 239 21847
rect 155 21687 239 21801
rect 155 21641 174 21687
rect 220 21641 239 21687
rect 155 21527 239 21641
rect 155 21481 174 21527
rect 220 21481 239 21527
rect 155 21367 239 21481
rect 155 21321 174 21367
rect 220 21321 239 21367
rect 155 21207 239 21321
rect 155 21161 174 21207
rect 220 21161 239 21207
rect 155 21047 239 21161
rect 155 21001 174 21047
rect 220 21001 239 21047
rect 155 20887 239 21001
rect 155 20841 174 20887
rect 220 20841 239 20887
rect 155 20727 239 20841
rect 155 20681 174 20727
rect 220 20681 239 20727
rect 155 20567 239 20681
rect 155 20521 174 20567
rect 220 20521 239 20567
rect 155 20407 239 20521
rect 155 20361 174 20407
rect 220 20361 239 20407
rect 155 20247 239 20361
rect 155 20201 174 20247
rect 220 20201 239 20247
rect 155 20087 239 20201
rect 155 20041 174 20087
rect 220 20041 239 20087
rect 155 19927 239 20041
rect 155 19881 174 19927
rect 220 19881 239 19927
rect 155 19767 239 19881
rect 155 19721 174 19767
rect 220 19721 239 19767
rect 155 19607 239 19721
rect 155 19561 174 19607
rect 220 19561 239 19607
rect 155 19447 239 19561
rect 155 19401 174 19447
rect 220 19401 239 19447
rect 155 19287 239 19401
rect 155 19241 174 19287
rect 220 19241 239 19287
rect 155 19127 239 19241
rect 155 19081 174 19127
rect 220 19081 239 19127
rect 155 18967 239 19081
rect 155 18921 174 18967
rect 220 18921 239 18967
rect 155 18807 239 18921
rect 155 18761 174 18807
rect 220 18761 239 18807
rect 155 18647 239 18761
rect 155 18601 174 18647
rect 220 18601 239 18647
rect 155 18487 239 18601
rect 155 18441 174 18487
rect 220 18441 239 18487
rect 155 18327 239 18441
rect 155 18281 174 18327
rect 220 18281 239 18327
rect 155 18167 239 18281
rect 155 18121 174 18167
rect 220 18121 239 18167
rect 155 18007 239 18121
rect 155 17961 174 18007
rect 220 17961 239 18007
rect 155 17847 239 17961
rect 155 17801 174 17847
rect 220 17801 239 17847
rect 155 17687 239 17801
rect 155 17641 174 17687
rect 220 17641 239 17687
rect 155 17527 239 17641
rect 155 17481 174 17527
rect 220 17481 239 17527
rect 155 17367 239 17481
rect 155 17321 174 17367
rect 220 17321 239 17367
rect 155 17207 239 17321
rect 155 17161 174 17207
rect 220 17161 239 17207
rect 155 17047 239 17161
rect 155 17001 174 17047
rect 220 17001 239 17047
rect 155 16887 239 17001
rect 155 16841 174 16887
rect 220 16841 239 16887
rect 155 16727 239 16841
rect 155 16681 174 16727
rect 220 16681 239 16727
rect 155 16567 239 16681
rect 155 16521 174 16567
rect 220 16521 239 16567
rect 155 16407 239 16521
rect 155 16361 174 16407
rect 220 16361 239 16407
rect 155 16247 239 16361
rect 155 16201 174 16247
rect 220 16201 239 16247
rect 155 16087 239 16201
rect 155 16041 174 16087
rect 220 16041 239 16087
rect 155 15927 239 16041
rect 155 15881 174 15927
rect 220 15881 239 15927
rect 155 15767 239 15881
rect 155 15721 174 15767
rect 220 15721 239 15767
rect 155 15607 239 15721
rect 155 15561 174 15607
rect 220 15561 239 15607
rect 155 15447 239 15561
rect 155 15401 174 15447
rect 220 15401 239 15447
rect 155 15287 239 15401
rect 155 15241 174 15287
rect 220 15241 239 15287
rect 155 15127 239 15241
rect 155 15081 174 15127
rect 220 15081 239 15127
rect 155 14967 239 15081
rect 155 14921 174 14967
rect 220 14921 239 14967
rect 155 14807 239 14921
rect 155 14761 174 14807
rect 220 14761 239 14807
rect 155 14647 239 14761
rect 155 14601 174 14647
rect 220 14601 239 14647
rect 155 14487 239 14601
rect 155 14441 174 14487
rect 220 14441 239 14487
rect 155 14327 239 14441
rect 155 14281 174 14327
rect 220 14281 239 14327
rect 155 14167 239 14281
rect 155 14121 174 14167
rect 220 14121 239 14167
rect 155 14007 239 14121
rect 155 13961 174 14007
rect 220 13961 239 14007
rect 155 13847 239 13961
rect 155 13801 174 13847
rect 220 13801 239 13847
rect 155 13687 239 13801
rect 155 13641 174 13687
rect 220 13641 239 13687
rect 155 13527 239 13641
rect 155 13481 174 13527
rect 220 13481 239 13527
rect 155 13386 239 13481
<< polycontact >>
rect 174 69641 220 69687
rect 174 69481 220 69527
rect 174 69321 220 69367
rect 174 69161 220 69207
rect 174 69001 220 69047
rect 174 68841 220 68887
rect 174 68681 220 68727
rect 174 68521 220 68567
rect 174 68361 220 68407
rect 174 68201 220 68247
rect 174 68041 220 68087
rect 174 67881 220 67927
rect 174 67721 220 67767
rect 174 67561 220 67607
rect 174 67401 220 67447
rect 174 67241 220 67287
rect 174 67081 220 67127
rect 174 66921 220 66967
rect 174 66761 220 66807
rect 174 66601 220 66647
rect 174 66441 220 66487
rect 174 66281 220 66327
rect 174 66121 220 66167
rect 174 65961 220 66007
rect 174 65801 220 65847
rect 174 65641 220 65687
rect 174 65481 220 65527
rect 174 65321 220 65367
rect 174 65161 220 65207
rect 174 65001 220 65047
rect 174 64841 220 64887
rect 174 64681 220 64727
rect 174 64521 220 64567
rect 174 64361 220 64407
rect 174 64201 220 64247
rect 174 64041 220 64087
rect 174 63881 220 63927
rect 174 63721 220 63767
rect 174 63561 220 63607
rect 174 63401 220 63447
rect 174 63241 220 63287
rect 174 63081 220 63127
rect 174 62921 220 62967
rect 174 62761 220 62807
rect 174 62601 220 62647
rect 174 62441 220 62487
rect 174 62281 220 62327
rect 174 62121 220 62167
rect 174 61961 220 62007
rect 174 61801 220 61847
rect 174 61641 220 61687
rect 174 61481 220 61527
rect 174 61321 220 61367
rect 174 61161 220 61207
rect 174 61001 220 61047
rect 174 60841 220 60887
rect 174 60681 220 60727
rect 174 60521 220 60567
rect 174 60361 220 60407
rect 174 60201 220 60247
rect 174 60041 220 60087
rect 174 59881 220 59927
rect 174 59721 220 59767
rect 174 59561 220 59607
rect 174 59401 220 59447
rect 174 59241 220 59287
rect 174 59081 220 59127
rect 174 58921 220 58967
rect 174 58761 220 58807
rect 174 58601 220 58647
rect 174 58441 220 58487
rect 174 58281 220 58327
rect 174 58121 220 58167
rect 174 57961 220 58007
rect 174 57801 220 57847
rect 174 57641 220 57687
rect 174 57481 220 57527
rect 174 57321 220 57367
rect 174 57161 220 57207
rect 174 57001 220 57047
rect 174 56841 220 56887
rect 174 56681 220 56727
rect 174 56521 220 56567
rect 174 56361 220 56407
rect 174 56201 220 56247
rect 174 56041 220 56087
rect 174 55881 220 55927
rect 174 55721 220 55767
rect 174 55561 220 55607
rect 174 55401 220 55447
rect 174 55241 220 55287
rect 174 55081 220 55127
rect 174 54921 220 54967
rect 174 54761 220 54807
rect 174 54601 220 54647
rect 174 54441 220 54487
rect 174 54281 220 54327
rect 174 54121 220 54167
rect 174 53961 220 54007
rect 174 53801 220 53847
rect 174 53641 220 53687
rect 174 53481 220 53527
rect 174 53321 220 53367
rect 174 53161 220 53207
rect 174 53001 220 53047
rect 174 52841 220 52887
rect 174 52681 220 52727
rect 174 52521 220 52567
rect 174 52361 220 52407
rect 174 52201 220 52247
rect 174 52041 220 52087
rect 174 51881 220 51927
rect 174 51721 220 51767
rect 174 51561 220 51607
rect 174 51401 220 51447
rect 174 51241 220 51287
rect 174 51081 220 51127
rect 174 50921 220 50967
rect 174 50761 220 50807
rect 174 50601 220 50647
rect 174 50441 220 50487
rect 174 50281 220 50327
rect 174 50121 220 50167
rect 174 49961 220 50007
rect 174 49801 220 49847
rect 174 49641 220 49687
rect 174 49481 220 49527
rect 174 49321 220 49367
rect 174 49161 220 49207
rect 174 49001 220 49047
rect 174 48841 220 48887
rect 174 48681 220 48727
rect 174 48521 220 48567
rect 174 48361 220 48407
rect 174 48201 220 48247
rect 174 48041 220 48087
rect 174 47881 220 47927
rect 174 47721 220 47767
rect 174 47561 220 47607
rect 174 47401 220 47447
rect 174 47241 220 47287
rect 174 47081 220 47127
rect 174 46921 220 46967
rect 174 46761 220 46807
rect 174 46601 220 46647
rect 174 46441 220 46487
rect 174 46281 220 46327
rect 174 46121 220 46167
rect 174 45961 220 46007
rect 174 45801 220 45847
rect 174 45641 220 45687
rect 174 45481 220 45527
rect 174 45321 220 45367
rect 174 45161 220 45207
rect 174 45001 220 45047
rect 174 44841 220 44887
rect 174 44681 220 44727
rect 174 44521 220 44567
rect 174 44361 220 44407
rect 174 44201 220 44247
rect 174 44041 220 44087
rect 174 43881 220 43927
rect 174 43721 220 43767
rect 174 43561 220 43607
rect 174 43401 220 43447
rect 174 43241 220 43287
rect 174 43081 220 43127
rect 174 42921 220 42967
rect 174 42761 220 42807
rect 174 42601 220 42647
rect 174 42441 220 42487
rect 174 42281 220 42327
rect 174 42121 220 42167
rect 174 41961 220 42007
rect 174 41801 220 41847
rect 174 41641 220 41687
rect 174 41481 220 41527
rect 174 41321 220 41367
rect 174 41161 220 41207
rect 174 41001 220 41047
rect 174 40841 220 40887
rect 174 40681 220 40727
rect 174 40521 220 40567
rect 174 40361 220 40407
rect 174 40201 220 40247
rect 174 40041 220 40087
rect 174 39881 220 39927
rect 174 39721 220 39767
rect 174 39561 220 39607
rect 174 39401 220 39447
rect 174 39241 220 39287
rect 174 39081 220 39127
rect 174 38921 220 38967
rect 174 38761 220 38807
rect 174 38601 220 38647
rect 174 38441 220 38487
rect 174 38281 220 38327
rect 174 38121 220 38167
rect 174 37961 220 38007
rect 174 37801 220 37847
rect 174 37641 220 37687
rect 174 37481 220 37527
rect 174 37321 220 37367
rect 174 37161 220 37207
rect 174 37001 220 37047
rect 174 36841 220 36887
rect 174 36681 220 36727
rect 174 36521 220 36567
rect 174 36361 220 36407
rect 174 36201 220 36247
rect 174 36041 220 36087
rect 174 35881 220 35927
rect 174 35721 220 35767
rect 174 35561 220 35607
rect 174 35401 220 35447
rect 174 35241 220 35287
rect 174 35081 220 35127
rect 174 34921 220 34967
rect 174 34761 220 34807
rect 174 34601 220 34647
rect 174 34441 220 34487
rect 174 34281 220 34327
rect 174 34121 220 34167
rect 174 33961 220 34007
rect 174 33801 220 33847
rect 174 33641 220 33687
rect 174 33481 220 33527
rect 174 33321 220 33367
rect 174 33161 220 33207
rect 174 33001 220 33047
rect 174 32841 220 32887
rect 174 32681 220 32727
rect 174 32521 220 32567
rect 174 32361 220 32407
rect 174 32201 220 32247
rect 174 32041 220 32087
rect 174 31881 220 31927
rect 174 31721 220 31767
rect 174 31561 220 31607
rect 174 31401 220 31447
rect 174 31241 220 31287
rect 174 31081 220 31127
rect 174 30921 220 30967
rect 174 30761 220 30807
rect 174 30601 220 30647
rect 174 30441 220 30487
rect 174 30281 220 30327
rect 174 30121 220 30167
rect 174 29961 220 30007
rect 174 29801 220 29847
rect 174 29641 220 29687
rect 174 29481 220 29527
rect 174 29321 220 29367
rect 174 29161 220 29207
rect 174 29001 220 29047
rect 174 28841 220 28887
rect 174 28681 220 28727
rect 174 28521 220 28567
rect 174 28361 220 28407
rect 174 28201 220 28247
rect 174 28041 220 28087
rect 174 27881 220 27927
rect 174 27721 220 27767
rect 174 27561 220 27607
rect 174 27401 220 27447
rect 174 27241 220 27287
rect 174 27081 220 27127
rect 174 26921 220 26967
rect 174 26761 220 26807
rect 174 26601 220 26647
rect 174 26441 220 26487
rect 174 26281 220 26327
rect 174 26121 220 26167
rect 174 25961 220 26007
rect 174 25801 220 25847
rect 174 25641 220 25687
rect 174 25481 220 25527
rect 174 25321 220 25367
rect 174 25161 220 25207
rect 174 25001 220 25047
rect 174 24841 220 24887
rect 174 24681 220 24727
rect 174 24521 220 24567
rect 174 24361 220 24407
rect 174 24201 220 24247
rect 174 24041 220 24087
rect 174 23881 220 23927
rect 174 23721 220 23767
rect 174 23561 220 23607
rect 174 23401 220 23447
rect 174 23241 220 23287
rect 174 23081 220 23127
rect 174 22921 220 22967
rect 174 22761 220 22807
rect 174 22601 220 22647
rect 174 22441 220 22487
rect 174 22281 220 22327
rect 174 22121 220 22167
rect 174 21961 220 22007
rect 174 21801 220 21847
rect 174 21641 220 21687
rect 174 21481 220 21527
rect 174 21321 220 21367
rect 174 21161 220 21207
rect 174 21001 220 21047
rect 174 20841 220 20887
rect 174 20681 220 20727
rect 174 20521 220 20567
rect 174 20361 220 20407
rect 174 20201 220 20247
rect 174 20041 220 20087
rect 174 19881 220 19927
rect 174 19721 220 19767
rect 174 19561 220 19607
rect 174 19401 220 19447
rect 174 19241 220 19287
rect 174 19081 220 19127
rect 174 18921 220 18967
rect 174 18761 220 18807
rect 174 18601 220 18647
rect 174 18441 220 18487
rect 174 18281 220 18327
rect 174 18121 220 18167
rect 174 17961 220 18007
rect 174 17801 220 17847
rect 174 17641 220 17687
rect 174 17481 220 17527
rect 174 17321 220 17367
rect 174 17161 220 17207
rect 174 17001 220 17047
rect 174 16841 220 16887
rect 174 16681 220 16727
rect 174 16521 220 16567
rect 174 16361 220 16407
rect 174 16201 220 16247
rect 174 16041 220 16087
rect 174 15881 220 15927
rect 174 15721 220 15767
rect 174 15561 220 15607
rect 174 15401 220 15447
rect 174 15241 220 15287
rect 174 15081 220 15127
rect 174 14921 220 14967
rect 174 14761 220 14807
rect 174 14601 220 14647
rect 174 14441 220 14487
rect 174 14281 220 14327
rect 174 14121 220 14167
rect 174 13961 220 14007
rect 174 13801 220 13847
rect 174 13641 220 13687
rect 174 13481 220 13527
<< metal1 >>
rect -32 69943 432 69957
rect -32 69871 130 69943
rect -32 69825 25 69871
rect 71 69825 130 69871
rect -32 69803 130 69825
rect 270 69871 432 69943
rect 270 69825 329 69871
rect 375 69825 432 69871
rect 270 69803 432 69825
rect -32 69789 432 69803
rect -32 69708 82 69789
rect -32 13356 25 69708
rect 71 69698 82 69708
rect 318 69708 432 69789
rect 318 69698 329 69708
rect 71 69687 329 69698
rect 71 69641 174 69687
rect 220 69641 329 69687
rect 71 69630 329 69641
rect 71 69538 82 69630
rect 318 69538 329 69630
rect 71 69527 329 69538
rect 71 69481 174 69527
rect 220 69481 329 69527
rect 71 69470 329 69481
rect 71 69378 82 69470
rect 318 69378 329 69470
rect 71 69367 329 69378
rect 71 69321 174 69367
rect 220 69321 329 69367
rect 71 69310 329 69321
rect 71 69218 82 69310
rect 318 69218 329 69310
rect 71 69207 329 69218
rect 71 69161 174 69207
rect 220 69161 329 69207
rect 71 69150 329 69161
rect 71 69058 82 69150
rect 318 69058 329 69150
rect 71 69047 329 69058
rect 71 69001 174 69047
rect 220 69001 329 69047
rect 71 68990 329 69001
rect 71 68898 82 68990
rect 318 68898 329 68990
rect 71 68887 329 68898
rect 71 68841 174 68887
rect 220 68841 329 68887
rect 71 68830 329 68841
rect 71 68738 82 68830
rect 318 68738 329 68830
rect 71 68727 329 68738
rect 71 68681 174 68727
rect 220 68681 329 68727
rect 71 68670 329 68681
rect 71 68578 82 68670
rect 318 68578 329 68670
rect 71 68567 329 68578
rect 71 68521 174 68567
rect 220 68521 329 68567
rect 71 68510 329 68521
rect 71 68418 82 68510
rect 318 68418 329 68510
rect 71 68407 329 68418
rect 71 68361 174 68407
rect 220 68361 329 68407
rect 71 68350 329 68361
rect 71 68258 82 68350
rect 318 68258 329 68350
rect 71 68247 329 68258
rect 71 68201 174 68247
rect 220 68201 329 68247
rect 71 68190 329 68201
rect 71 68098 82 68190
rect 318 68098 329 68190
rect 71 68087 329 68098
rect 71 68041 174 68087
rect 220 68041 329 68087
rect 71 68030 329 68041
rect 71 67938 82 68030
rect 318 67938 329 68030
rect 71 67927 329 67938
rect 71 67881 174 67927
rect 220 67881 329 67927
rect 71 67870 329 67881
rect 71 67778 82 67870
rect 318 67778 329 67870
rect 71 67767 329 67778
rect 71 67721 174 67767
rect 220 67721 329 67767
rect 71 67710 329 67721
rect 71 67618 82 67710
rect 318 67618 329 67710
rect 71 67607 329 67618
rect 71 67561 174 67607
rect 220 67561 329 67607
rect 71 67550 329 67561
rect 71 67458 82 67550
rect 318 67458 329 67550
rect 71 67447 329 67458
rect 71 67401 174 67447
rect 220 67401 329 67447
rect 71 67390 329 67401
rect 71 67298 82 67390
rect 318 67298 329 67390
rect 71 67287 329 67298
rect 71 67241 174 67287
rect 220 67241 329 67287
rect 71 67230 329 67241
rect 71 67138 82 67230
rect 318 67138 329 67230
rect 71 67127 329 67138
rect 71 67081 174 67127
rect 220 67081 329 67127
rect 71 67070 329 67081
rect 71 66978 82 67070
rect 318 66978 329 67070
rect 71 66967 329 66978
rect 71 66921 174 66967
rect 220 66921 329 66967
rect 71 66910 329 66921
rect 71 66818 82 66910
rect 318 66818 329 66910
rect 71 66807 329 66818
rect 71 66761 174 66807
rect 220 66761 329 66807
rect 71 66750 329 66761
rect 71 66658 82 66750
rect 318 66658 329 66750
rect 71 66647 329 66658
rect 71 66601 174 66647
rect 220 66601 329 66647
rect 71 66590 329 66601
rect 71 66498 82 66590
rect 318 66498 329 66590
rect 71 66487 329 66498
rect 71 66441 174 66487
rect 220 66441 329 66487
rect 71 66430 329 66441
rect 71 66338 82 66430
rect 318 66338 329 66430
rect 71 66327 329 66338
rect 71 66281 174 66327
rect 220 66281 329 66327
rect 71 66270 329 66281
rect 71 66178 82 66270
rect 318 66178 329 66270
rect 71 66167 329 66178
rect 71 66121 174 66167
rect 220 66121 329 66167
rect 71 66110 329 66121
rect 71 66018 82 66110
rect 318 66018 329 66110
rect 71 66007 329 66018
rect 71 65961 174 66007
rect 220 65961 329 66007
rect 71 65950 329 65961
rect 71 65858 82 65950
rect 318 65858 329 65950
rect 71 65847 329 65858
rect 71 65801 174 65847
rect 220 65801 329 65847
rect 71 65790 329 65801
rect 71 65698 82 65790
rect 318 65698 329 65790
rect 71 65687 329 65698
rect 71 65641 174 65687
rect 220 65641 329 65687
rect 71 65630 329 65641
rect 71 65538 82 65630
rect 318 65538 329 65630
rect 71 65527 329 65538
rect 71 65481 174 65527
rect 220 65481 329 65527
rect 71 65470 329 65481
rect 71 65378 82 65470
rect 318 65378 329 65470
rect 71 65367 329 65378
rect 71 65321 174 65367
rect 220 65321 329 65367
rect 71 65310 329 65321
rect 71 65218 82 65310
rect 318 65218 329 65310
rect 71 65207 329 65218
rect 71 65161 174 65207
rect 220 65161 329 65207
rect 71 65150 329 65161
rect 71 65058 82 65150
rect 318 65058 329 65150
rect 71 65047 329 65058
rect 71 65001 174 65047
rect 220 65001 329 65047
rect 71 64942 329 65001
rect 71 64890 130 64942
rect 286 64890 329 64942
rect 71 64887 329 64890
rect 71 64841 174 64887
rect 220 64841 329 64887
rect 71 64830 329 64841
rect 71 64778 130 64830
rect 286 64778 329 64830
rect 71 64727 329 64778
rect 71 64718 174 64727
rect 220 64718 329 64727
rect 71 64666 130 64718
rect 286 64666 329 64718
rect 71 64606 329 64666
rect 71 64554 130 64606
rect 286 64554 329 64606
rect 71 64521 174 64554
rect 220 64521 329 64554
rect 71 64494 329 64521
rect 71 64442 130 64494
rect 286 64442 329 64494
rect 71 64407 329 64442
rect 71 64382 174 64407
rect 220 64382 329 64407
rect 71 64330 130 64382
rect 286 64330 329 64382
rect 71 64270 329 64330
rect 71 64218 130 64270
rect 286 64218 329 64270
rect 71 64201 174 64218
rect 220 64201 329 64218
rect 71 64158 329 64201
rect 71 64106 130 64158
rect 286 64106 329 64158
rect 71 64087 329 64106
rect 71 64046 174 64087
rect 220 64046 329 64087
rect 71 63994 130 64046
rect 286 63994 329 64046
rect 71 63934 329 63994
rect 71 63882 130 63934
rect 286 63882 329 63934
rect 71 63881 174 63882
rect 220 63881 329 63882
rect 71 63822 329 63881
rect 71 63770 130 63822
rect 286 63770 329 63822
rect 71 63767 329 63770
rect 71 63721 174 63767
rect 220 63721 329 63767
rect 71 63710 329 63721
rect 71 63658 130 63710
rect 286 63658 329 63710
rect 71 63607 329 63658
rect 71 63561 174 63607
rect 220 63561 329 63607
rect 71 63550 329 63561
rect 71 63458 82 63550
rect 318 63458 329 63550
rect 71 63447 329 63458
rect 71 63401 174 63447
rect 220 63401 329 63447
rect 71 63390 329 63401
rect 71 63298 82 63390
rect 318 63298 329 63390
rect 71 63287 329 63298
rect 71 63241 174 63287
rect 220 63241 329 63287
rect 71 63230 329 63241
rect 71 63138 82 63230
rect 318 63138 329 63230
rect 71 63127 329 63138
rect 71 63081 174 63127
rect 220 63081 329 63127
rect 71 63070 329 63081
rect 71 62978 82 63070
rect 318 62978 329 63070
rect 71 62967 329 62978
rect 71 62921 174 62967
rect 220 62921 329 62967
rect 71 62910 329 62921
rect 71 62818 82 62910
rect 318 62818 329 62910
rect 71 62807 329 62818
rect 71 62761 174 62807
rect 220 62761 329 62807
rect 71 62750 329 62761
rect 71 62658 82 62750
rect 318 62658 329 62750
rect 71 62647 329 62658
rect 71 62601 174 62647
rect 220 62601 329 62647
rect 71 62590 329 62601
rect 71 62498 82 62590
rect 318 62498 329 62590
rect 71 62487 329 62498
rect 71 62441 174 62487
rect 220 62441 329 62487
rect 71 62430 329 62441
rect 71 62338 82 62430
rect 318 62338 329 62430
rect 71 62327 329 62338
rect 71 62281 174 62327
rect 220 62281 329 62327
rect 71 62270 329 62281
rect 71 62178 82 62270
rect 318 62178 329 62270
rect 71 62167 329 62178
rect 71 62121 174 62167
rect 220 62121 329 62167
rect 71 62110 329 62121
rect 71 62018 82 62110
rect 318 62018 329 62110
rect 71 62007 329 62018
rect 71 61961 174 62007
rect 220 61961 329 62007
rect 71 61950 329 61961
rect 71 61858 82 61950
rect 318 61858 329 61950
rect 71 61847 329 61858
rect 71 61801 174 61847
rect 220 61801 329 61847
rect 71 61790 329 61801
rect 71 61698 82 61790
rect 318 61698 329 61790
rect 71 61687 329 61698
rect 71 61641 174 61687
rect 220 61641 329 61687
rect 71 61630 329 61641
rect 71 61538 82 61630
rect 318 61538 329 61630
rect 71 61527 329 61538
rect 71 61481 174 61527
rect 220 61481 329 61527
rect 71 61470 329 61481
rect 71 61378 82 61470
rect 318 61378 329 61470
rect 71 61367 329 61378
rect 71 61321 174 61367
rect 220 61321 329 61367
rect 71 61310 329 61321
rect 71 61218 82 61310
rect 318 61218 329 61310
rect 71 61207 329 61218
rect 71 61161 174 61207
rect 220 61161 329 61207
rect 71 61150 329 61161
rect 71 61058 82 61150
rect 318 61058 329 61150
rect 71 61047 329 61058
rect 71 61001 174 61047
rect 220 61001 329 61047
rect 71 60990 329 61001
rect 71 60898 82 60990
rect 318 60898 329 60990
rect 71 60887 329 60898
rect 71 60841 174 60887
rect 220 60841 329 60887
rect 71 60830 329 60841
rect 71 60738 82 60830
rect 318 60738 329 60830
rect 71 60727 329 60738
rect 71 60681 174 60727
rect 220 60681 329 60727
rect 71 60670 329 60681
rect 71 60578 82 60670
rect 318 60578 329 60670
rect 71 60567 329 60578
rect 71 60521 174 60567
rect 220 60521 329 60567
rect 71 60510 329 60521
rect 71 60418 82 60510
rect 318 60418 329 60510
rect 71 60407 329 60418
rect 71 60361 174 60407
rect 220 60361 329 60407
rect 71 60350 329 60361
rect 71 60258 82 60350
rect 318 60258 329 60350
rect 71 60247 329 60258
rect 71 60201 174 60247
rect 220 60201 329 60247
rect 71 60190 329 60201
rect 71 60098 82 60190
rect 318 60098 329 60190
rect 71 60087 329 60098
rect 71 60041 174 60087
rect 220 60041 329 60087
rect 71 60030 329 60041
rect 71 59938 82 60030
rect 318 59938 329 60030
rect 71 59927 329 59938
rect 71 59881 174 59927
rect 220 59881 329 59927
rect 71 59870 329 59881
rect 71 59778 82 59870
rect 318 59778 329 59870
rect 71 59767 329 59778
rect 71 59721 174 59767
rect 220 59721 329 59767
rect 71 59710 329 59721
rect 71 59618 82 59710
rect 318 59618 329 59710
rect 71 59607 329 59618
rect 71 59561 174 59607
rect 220 59561 329 59607
rect 71 59550 329 59561
rect 71 59458 82 59550
rect 318 59458 329 59550
rect 71 59447 329 59458
rect 71 59401 174 59447
rect 220 59401 329 59447
rect 71 59390 329 59401
rect 71 59298 82 59390
rect 318 59298 329 59390
rect 71 59287 329 59298
rect 71 59241 174 59287
rect 220 59241 329 59287
rect 71 59230 329 59241
rect 71 59138 82 59230
rect 318 59138 329 59230
rect 71 59127 329 59138
rect 71 59081 174 59127
rect 220 59081 329 59127
rect 71 59070 329 59081
rect 71 58978 82 59070
rect 318 58978 329 59070
rect 71 58967 329 58978
rect 71 58921 174 58967
rect 220 58921 329 58967
rect 71 58910 329 58921
rect 71 58818 82 58910
rect 318 58818 329 58910
rect 71 58807 329 58818
rect 71 58761 174 58807
rect 220 58761 329 58807
rect 71 58750 329 58761
rect 71 58658 82 58750
rect 318 58658 329 58750
rect 71 58647 329 58658
rect 71 58601 174 58647
rect 220 58601 329 58647
rect 71 58590 329 58601
rect 71 58498 82 58590
rect 318 58498 329 58590
rect 71 58487 329 58498
rect 71 58441 174 58487
rect 220 58441 329 58487
rect 71 58430 329 58441
rect 71 58338 82 58430
rect 318 58338 329 58430
rect 71 58327 329 58338
rect 71 58281 174 58327
rect 220 58281 329 58327
rect 71 58270 329 58281
rect 71 58178 82 58270
rect 318 58178 329 58270
rect 71 58167 329 58178
rect 71 58121 174 58167
rect 220 58121 329 58167
rect 71 58110 329 58121
rect 71 58018 82 58110
rect 318 58018 329 58110
rect 71 58007 329 58018
rect 71 57961 174 58007
rect 220 57961 329 58007
rect 71 57950 329 57961
rect 71 57858 82 57950
rect 318 57858 329 57950
rect 71 57847 329 57858
rect 71 57801 174 57847
rect 220 57801 329 57847
rect 71 57790 329 57801
rect 71 57698 82 57790
rect 318 57698 329 57790
rect 71 57687 329 57698
rect 71 57641 174 57687
rect 220 57641 329 57687
rect 71 57630 329 57641
rect 71 57538 82 57630
rect 318 57538 329 57630
rect 71 57527 329 57538
rect 71 57481 174 57527
rect 220 57481 329 57527
rect 71 57470 329 57481
rect 71 57378 82 57470
rect 318 57378 329 57470
rect 71 57367 329 57378
rect 71 57321 174 57367
rect 220 57321 329 57367
rect 71 57310 329 57321
rect 71 57218 82 57310
rect 318 57218 329 57310
rect 71 57207 329 57218
rect 71 57161 174 57207
rect 220 57161 329 57207
rect 71 57150 329 57161
rect 71 57058 82 57150
rect 318 57058 329 57150
rect 71 57047 329 57058
rect 71 57001 174 57047
rect 220 57001 329 57047
rect 71 56990 329 57001
rect 71 56898 82 56990
rect 318 56898 329 56990
rect 71 56887 329 56898
rect 71 56841 174 56887
rect 220 56841 329 56887
rect 71 56830 329 56841
rect 71 56738 82 56830
rect 318 56738 329 56830
rect 71 56727 329 56738
rect 71 56681 174 56727
rect 220 56681 329 56727
rect 71 56670 329 56681
rect 71 56578 82 56670
rect 318 56578 329 56670
rect 71 56567 329 56578
rect 71 56521 174 56567
rect 220 56521 329 56567
rect 71 56510 329 56521
rect 71 56418 82 56510
rect 318 56418 329 56510
rect 71 56407 329 56418
rect 71 56361 174 56407
rect 220 56361 329 56407
rect 71 56350 329 56361
rect 71 56258 82 56350
rect 318 56258 329 56350
rect 71 56247 329 56258
rect 71 56201 174 56247
rect 220 56201 329 56247
rect 71 56190 329 56201
rect 71 56098 82 56190
rect 318 56098 329 56190
rect 71 56087 329 56098
rect 71 56041 174 56087
rect 220 56041 329 56087
rect 71 56030 329 56041
rect 71 55938 82 56030
rect 318 55938 329 56030
rect 71 55927 329 55938
rect 71 55881 174 55927
rect 220 55881 329 55927
rect 71 55870 329 55881
rect 71 55778 82 55870
rect 318 55778 329 55870
rect 71 55767 329 55778
rect 71 55721 174 55767
rect 220 55721 329 55767
rect 71 55710 329 55721
rect 71 55618 82 55710
rect 318 55618 329 55710
rect 71 55607 329 55618
rect 71 55561 174 55607
rect 220 55561 329 55607
rect 71 55550 329 55561
rect 71 55458 82 55550
rect 318 55458 329 55550
rect 71 55447 329 55458
rect 71 55401 174 55447
rect 220 55401 329 55447
rect 71 55390 329 55401
rect 71 55298 82 55390
rect 318 55298 329 55390
rect 71 55287 329 55298
rect 71 55241 174 55287
rect 220 55241 329 55287
rect 71 55230 329 55241
rect 71 55138 82 55230
rect 318 55138 329 55230
rect 71 55127 329 55138
rect 71 55081 174 55127
rect 220 55081 329 55127
rect 71 55070 329 55081
rect 71 54978 82 55070
rect 318 54978 329 55070
rect 71 54967 329 54978
rect 71 54921 174 54967
rect 220 54921 329 54967
rect 71 54910 329 54921
rect 71 54818 82 54910
rect 318 54818 329 54910
rect 71 54807 329 54818
rect 71 54761 174 54807
rect 220 54761 329 54807
rect 71 54750 329 54761
rect 71 54658 82 54750
rect 318 54658 329 54750
rect 71 54647 329 54658
rect 71 54601 174 54647
rect 220 54601 329 54647
rect 71 54590 329 54601
rect 71 54498 82 54590
rect 318 54498 329 54590
rect 71 54487 329 54498
rect 71 54441 174 54487
rect 220 54441 329 54487
rect 71 54430 329 54441
rect 71 54338 82 54430
rect 318 54338 329 54430
rect 71 54327 329 54338
rect 71 54281 174 54327
rect 220 54281 329 54327
rect 71 54270 329 54281
rect 71 54178 82 54270
rect 318 54178 329 54270
rect 71 54167 329 54178
rect 71 54121 174 54167
rect 220 54121 329 54167
rect 71 54110 329 54121
rect 71 54018 82 54110
rect 318 54018 329 54110
rect 71 54007 329 54018
rect 71 53961 174 54007
rect 220 53961 329 54007
rect 71 53950 329 53961
rect 71 53858 82 53950
rect 318 53858 329 53950
rect 71 53847 329 53858
rect 71 53801 174 53847
rect 220 53801 329 53847
rect 71 53790 329 53801
rect 71 53698 82 53790
rect 318 53698 329 53790
rect 71 53687 329 53698
rect 71 53641 174 53687
rect 220 53641 329 53687
rect 71 53630 329 53641
rect 71 53538 82 53630
rect 318 53538 329 53630
rect 71 53527 329 53538
rect 71 53481 174 53527
rect 220 53481 329 53527
rect 71 53470 329 53481
rect 71 53378 82 53470
rect 318 53378 329 53470
rect 71 53367 329 53378
rect 71 53321 174 53367
rect 220 53321 329 53367
rect 71 53310 329 53321
rect 71 53218 82 53310
rect 318 53218 329 53310
rect 71 53207 329 53218
rect 71 53161 174 53207
rect 220 53161 329 53207
rect 71 53150 329 53161
rect 71 53058 82 53150
rect 318 53058 329 53150
rect 71 53047 329 53058
rect 71 53001 174 53047
rect 220 53001 329 53047
rect 71 52990 329 53001
rect 71 52898 82 52990
rect 318 52898 329 52990
rect 71 52887 329 52898
rect 71 52841 174 52887
rect 220 52841 329 52887
rect 71 52830 329 52841
rect 71 52738 82 52830
rect 318 52738 329 52830
rect 71 52727 329 52738
rect 71 52681 174 52727
rect 220 52681 329 52727
rect 71 52670 329 52681
rect 71 52578 82 52670
rect 318 52578 329 52670
rect 71 52567 329 52578
rect 71 52521 174 52567
rect 220 52521 329 52567
rect 71 52510 329 52521
rect 71 52418 82 52510
rect 318 52418 329 52510
rect 71 52407 329 52418
rect 71 52361 174 52407
rect 220 52361 329 52407
rect 71 52350 329 52361
rect 71 52258 82 52350
rect 318 52258 329 52350
rect 71 52247 329 52258
rect 71 52201 174 52247
rect 220 52201 329 52247
rect 71 52190 329 52201
rect 71 52098 82 52190
rect 318 52098 329 52190
rect 71 52087 329 52098
rect 71 52041 174 52087
rect 220 52041 329 52087
rect 71 52030 329 52041
rect 71 51938 82 52030
rect 318 51938 329 52030
rect 71 51927 329 51938
rect 71 51881 174 51927
rect 220 51881 329 51927
rect 71 51870 329 51881
rect 71 51778 82 51870
rect 318 51778 329 51870
rect 71 51767 329 51778
rect 71 51721 174 51767
rect 220 51721 329 51767
rect 71 51710 329 51721
rect 71 51618 82 51710
rect 318 51618 329 51710
rect 71 51607 329 51618
rect 71 51561 174 51607
rect 220 51561 329 51607
rect 71 51550 329 51561
rect 71 51458 82 51550
rect 318 51458 329 51550
rect 71 51447 329 51458
rect 71 51401 174 51447
rect 220 51401 329 51447
rect 71 51390 329 51401
rect 71 51298 82 51390
rect 318 51298 329 51390
rect 71 51287 329 51298
rect 71 51241 174 51287
rect 220 51241 329 51287
rect 71 51230 329 51241
rect 71 51138 82 51230
rect 318 51138 329 51230
rect 71 51127 329 51138
rect 71 51081 174 51127
rect 220 51081 329 51127
rect 71 51070 329 51081
rect 71 50978 82 51070
rect 318 50978 329 51070
rect 71 50967 329 50978
rect 71 50921 174 50967
rect 220 50921 329 50967
rect 71 50910 329 50921
rect 71 50818 82 50910
rect 318 50818 329 50910
rect 71 50807 329 50818
rect 71 50761 174 50807
rect 220 50761 329 50807
rect 71 50750 329 50761
rect 71 50658 82 50750
rect 318 50658 329 50750
rect 71 50647 329 50658
rect 71 50601 174 50647
rect 220 50601 329 50647
rect 71 50536 329 50601
rect 71 50484 127 50536
rect 179 50487 239 50536
rect 220 50484 239 50487
rect 291 50484 329 50536
rect 71 50441 174 50484
rect 220 50441 329 50484
rect 71 50424 329 50441
rect 71 50372 127 50424
rect 179 50372 239 50424
rect 291 50372 329 50424
rect 71 50327 329 50372
rect 71 50312 174 50327
rect 220 50312 329 50327
rect 71 50260 127 50312
rect 220 50281 239 50312
rect 179 50260 239 50281
rect 291 50260 329 50312
rect 71 50200 329 50260
rect 71 50148 127 50200
rect 179 50167 239 50200
rect 220 50148 239 50167
rect 291 50148 329 50200
rect 71 50121 174 50148
rect 220 50121 329 50148
rect 71 50088 329 50121
rect 71 50036 127 50088
rect 179 50036 239 50088
rect 291 50036 329 50088
rect 71 50007 329 50036
rect 71 49976 174 50007
rect 220 49976 329 50007
rect 71 49924 127 49976
rect 220 49961 239 49976
rect 179 49924 239 49961
rect 291 49924 329 49976
rect 71 49864 329 49924
rect 71 49812 127 49864
rect 179 49847 239 49864
rect 220 49812 239 49847
rect 291 49812 329 49864
rect 71 49801 174 49812
rect 220 49801 329 49812
rect 71 49752 329 49801
rect 71 49700 127 49752
rect 179 49700 239 49752
rect 291 49700 329 49752
rect 71 49687 329 49700
rect 71 49641 174 49687
rect 220 49641 329 49687
rect 71 49640 329 49641
rect 71 49588 127 49640
rect 179 49588 239 49640
rect 291 49588 329 49640
rect 71 49528 329 49588
rect 71 49476 127 49528
rect 179 49527 239 49528
rect 220 49481 239 49527
rect 179 49476 239 49481
rect 291 49476 329 49528
rect 71 49416 329 49476
rect 71 49364 127 49416
rect 179 49367 239 49416
rect 220 49364 239 49367
rect 291 49364 329 49416
rect 71 49321 174 49364
rect 220 49321 329 49364
rect 71 49304 329 49321
rect 71 49252 127 49304
rect 179 49252 239 49304
rect 291 49252 329 49304
rect 71 49207 329 49252
rect 71 49161 174 49207
rect 220 49161 329 49207
rect 71 49150 329 49161
rect 71 49058 82 49150
rect 318 49058 329 49150
rect 71 49047 329 49058
rect 71 49001 174 49047
rect 220 49001 329 49047
rect 71 48990 329 49001
rect 71 48898 82 48990
rect 318 48898 329 48990
rect 71 48887 329 48898
rect 71 48841 174 48887
rect 220 48841 329 48887
rect 71 48830 329 48841
rect 71 48738 82 48830
rect 318 48738 329 48830
rect 71 48727 329 48738
rect 71 48681 174 48727
rect 220 48681 329 48727
rect 71 48670 329 48681
rect 71 48578 82 48670
rect 318 48578 329 48670
rect 71 48567 329 48578
rect 71 48521 174 48567
rect 220 48521 329 48567
rect 71 48510 329 48521
rect 71 48418 82 48510
rect 318 48418 329 48510
rect 71 48407 329 48418
rect 71 48361 174 48407
rect 220 48361 329 48407
rect 71 48350 329 48361
rect 71 48258 82 48350
rect 318 48258 329 48350
rect 71 48247 329 48258
rect 71 48201 174 48247
rect 220 48201 329 48247
rect 71 48190 329 48201
rect 71 48098 82 48190
rect 318 48098 329 48190
rect 71 48087 329 48098
rect 71 48041 174 48087
rect 220 48041 329 48087
rect 71 48030 329 48041
rect 71 47938 82 48030
rect 318 47938 329 48030
rect 71 47927 329 47938
rect 71 47881 174 47927
rect 220 47881 329 47927
rect 71 47870 329 47881
rect 71 47778 82 47870
rect 318 47778 329 47870
rect 71 47767 329 47778
rect 71 47721 174 47767
rect 220 47721 329 47767
rect 71 47710 329 47721
rect 71 47618 82 47710
rect 318 47618 329 47710
rect 71 47607 329 47618
rect 71 47561 174 47607
rect 220 47561 329 47607
rect 71 47550 329 47561
rect 71 47458 82 47550
rect 318 47458 329 47550
rect 71 47447 329 47458
rect 71 47401 174 47447
rect 220 47401 329 47447
rect 71 47390 329 47401
rect 71 47298 82 47390
rect 318 47298 329 47390
rect 71 47287 329 47298
rect 71 47241 174 47287
rect 220 47241 329 47287
rect 71 47230 329 47241
rect 71 47138 82 47230
rect 318 47138 329 47230
rect 71 47127 329 47138
rect 71 47081 174 47127
rect 220 47081 329 47127
rect 71 47070 329 47081
rect 71 46978 82 47070
rect 318 46978 329 47070
rect 71 46967 329 46978
rect 71 46921 174 46967
rect 220 46921 329 46967
rect 71 46910 329 46921
rect 71 46818 82 46910
rect 318 46818 329 46910
rect 71 46807 329 46818
rect 71 46761 174 46807
rect 220 46761 329 46807
rect 71 46750 329 46761
rect 71 46658 82 46750
rect 318 46658 329 46750
rect 71 46647 329 46658
rect 71 46601 174 46647
rect 220 46601 329 46647
rect 71 46590 329 46601
rect 71 46498 82 46590
rect 318 46498 329 46590
rect 71 46487 329 46498
rect 71 46441 174 46487
rect 220 46441 329 46487
rect 71 46430 329 46441
rect 71 46338 82 46430
rect 318 46338 329 46430
rect 71 46327 329 46338
rect 71 46281 174 46327
rect 220 46281 329 46327
rect 71 46270 329 46281
rect 71 46178 82 46270
rect 318 46178 329 46270
rect 71 46167 329 46178
rect 71 46121 174 46167
rect 220 46121 329 46167
rect 71 46110 329 46121
rect 71 46018 82 46110
rect 318 46018 329 46110
rect 71 46007 329 46018
rect 71 45961 174 46007
rect 220 45961 329 46007
rect 71 45950 329 45961
rect 71 45858 82 45950
rect 318 45858 329 45950
rect 71 45847 329 45858
rect 71 45801 174 45847
rect 220 45801 329 45847
rect 71 45790 329 45801
rect 71 45698 82 45790
rect 318 45698 329 45790
rect 71 45687 329 45698
rect 71 45641 174 45687
rect 220 45641 329 45687
rect 71 45630 329 45641
rect 71 45538 82 45630
rect 318 45538 329 45630
rect 71 45527 329 45538
rect 71 45481 174 45527
rect 220 45481 329 45527
rect 71 45470 329 45481
rect 71 45378 82 45470
rect 318 45378 329 45470
rect 71 45367 329 45378
rect 71 45321 174 45367
rect 220 45321 329 45367
rect 71 45310 329 45321
rect 71 45218 82 45310
rect 318 45218 329 45310
rect 71 45207 329 45218
rect 71 45161 174 45207
rect 220 45161 329 45207
rect 71 45150 329 45161
rect 71 45058 82 45150
rect 318 45058 329 45150
rect 71 45047 329 45058
rect 71 45001 174 45047
rect 220 45001 329 45047
rect 71 44990 329 45001
rect 71 44898 82 44990
rect 318 44898 329 44990
rect 71 44887 329 44898
rect 71 44841 174 44887
rect 220 44841 329 44887
rect 71 44830 329 44841
rect 71 44738 82 44830
rect 318 44738 329 44830
rect 71 44727 329 44738
rect 71 44681 174 44727
rect 220 44681 329 44727
rect 71 44670 329 44681
rect 71 44578 82 44670
rect 318 44578 329 44670
rect 71 44567 329 44578
rect 71 44521 174 44567
rect 220 44521 329 44567
rect 71 44510 329 44521
rect 71 44418 82 44510
rect 318 44418 329 44510
rect 71 44407 329 44418
rect 71 44361 174 44407
rect 220 44361 329 44407
rect 71 44350 329 44361
rect 71 44258 82 44350
rect 318 44258 329 44350
rect 71 44247 329 44258
rect 71 44201 174 44247
rect 220 44201 329 44247
rect 71 44190 329 44201
rect 71 44098 82 44190
rect 318 44098 329 44190
rect 71 44087 329 44098
rect 71 44041 174 44087
rect 220 44041 329 44087
rect 71 44030 329 44041
rect 71 43938 82 44030
rect 318 43938 329 44030
rect 71 43927 329 43938
rect 71 43881 174 43927
rect 220 43881 329 43927
rect 71 43870 329 43881
rect 71 43778 82 43870
rect 318 43778 329 43870
rect 71 43767 329 43778
rect 71 43721 174 43767
rect 220 43721 329 43767
rect 71 43710 329 43721
rect 71 43618 82 43710
rect 318 43618 329 43710
rect 71 43607 329 43618
rect 71 43561 174 43607
rect 220 43561 329 43607
rect 71 43550 329 43561
rect 71 43458 82 43550
rect 318 43458 329 43550
rect 71 43447 329 43458
rect 71 43401 174 43447
rect 220 43401 329 43447
rect 71 43390 329 43401
rect 71 43298 82 43390
rect 318 43298 329 43390
rect 71 43287 329 43298
rect 71 43241 174 43287
rect 220 43241 329 43287
rect 71 43230 329 43241
rect 71 43138 82 43230
rect 318 43138 329 43230
rect 71 43127 329 43138
rect 71 43081 174 43127
rect 220 43081 329 43127
rect 71 43070 329 43081
rect 71 42978 82 43070
rect 318 42978 329 43070
rect 71 42967 329 42978
rect 71 42921 174 42967
rect 220 42921 329 42967
rect 71 42910 329 42921
rect 71 42818 82 42910
rect 318 42818 329 42910
rect 71 42807 329 42818
rect 71 42761 174 42807
rect 220 42761 329 42807
rect 71 42750 329 42761
rect 71 42658 82 42750
rect 318 42658 329 42750
rect 71 42647 329 42658
rect 71 42601 174 42647
rect 220 42601 329 42647
rect 71 42590 329 42601
rect 71 42498 82 42590
rect 318 42498 329 42590
rect 71 42487 329 42498
rect 71 42441 174 42487
rect 220 42441 329 42487
rect 71 42430 329 42441
rect 71 42338 82 42430
rect 318 42338 329 42430
rect 71 42327 329 42338
rect 71 42281 174 42327
rect 220 42281 329 42327
rect 71 42270 329 42281
rect 71 42178 82 42270
rect 318 42178 329 42270
rect 71 42167 329 42178
rect 71 42121 174 42167
rect 220 42121 329 42167
rect 71 42110 329 42121
rect 71 42018 82 42110
rect 318 42018 329 42110
rect 71 42007 329 42018
rect 71 41961 174 42007
rect 220 41961 329 42007
rect 71 41950 329 41961
rect 71 41858 82 41950
rect 318 41858 329 41950
rect 71 41847 329 41858
rect 71 41801 174 41847
rect 220 41801 329 41847
rect 71 41790 329 41801
rect 71 41698 82 41790
rect 318 41698 329 41790
rect 71 41687 329 41698
rect 71 41641 174 41687
rect 220 41641 329 41687
rect 71 41630 329 41641
rect 71 41538 82 41630
rect 318 41538 329 41630
rect 71 41527 329 41538
rect 71 41481 174 41527
rect 220 41481 329 41527
rect 71 41470 329 41481
rect 71 41378 82 41470
rect 318 41378 329 41470
rect 71 41367 329 41378
rect 71 41321 174 41367
rect 220 41321 329 41367
rect 71 41310 329 41321
rect 71 41218 82 41310
rect 318 41218 329 41310
rect 71 41207 329 41218
rect 71 41161 174 41207
rect 220 41161 329 41207
rect 71 41150 329 41161
rect 71 41058 82 41150
rect 318 41058 329 41150
rect 71 41047 329 41058
rect 71 41001 174 41047
rect 220 41001 329 41047
rect 71 40990 329 41001
rect 71 40898 82 40990
rect 318 40898 329 40990
rect 71 40887 329 40898
rect 71 40841 174 40887
rect 220 40841 329 40887
rect 71 40830 329 40841
rect 71 40738 82 40830
rect 318 40738 329 40830
rect 71 40727 329 40738
rect 71 40681 174 40727
rect 220 40681 329 40727
rect 71 40670 329 40681
rect 71 40578 82 40670
rect 318 40578 329 40670
rect 71 40567 329 40578
rect 71 40521 174 40567
rect 220 40521 329 40567
rect 71 40510 329 40521
rect 71 40418 82 40510
rect 318 40418 329 40510
rect 71 40407 329 40418
rect 71 40361 174 40407
rect 220 40361 329 40407
rect 71 40350 329 40361
rect 71 40258 82 40350
rect 318 40258 329 40350
rect 71 40247 329 40258
rect 71 40201 174 40247
rect 220 40201 329 40247
rect 71 40190 329 40201
rect 71 40098 82 40190
rect 318 40098 329 40190
rect 71 40087 329 40098
rect 71 40041 174 40087
rect 220 40041 329 40087
rect 71 40030 329 40041
rect 71 39938 82 40030
rect 318 39938 329 40030
rect 71 39927 329 39938
rect 71 39881 174 39927
rect 220 39881 329 39927
rect 71 39870 329 39881
rect 71 39778 82 39870
rect 318 39778 329 39870
rect 71 39767 329 39778
rect 71 39721 174 39767
rect 220 39721 329 39767
rect 71 39710 329 39721
rect 71 39618 82 39710
rect 318 39618 329 39710
rect 71 39607 329 39618
rect 71 39561 174 39607
rect 220 39561 329 39607
rect 71 39550 329 39561
rect 71 39458 82 39550
rect 318 39458 329 39550
rect 71 39447 329 39458
rect 71 39401 174 39447
rect 220 39401 329 39447
rect 71 39390 329 39401
rect 71 39298 82 39390
rect 318 39298 329 39390
rect 71 39287 329 39298
rect 71 39241 174 39287
rect 220 39241 329 39287
rect 71 39230 329 39241
rect 71 39138 82 39230
rect 318 39138 329 39230
rect 71 39127 329 39138
rect 71 39081 174 39127
rect 220 39081 329 39127
rect 71 39070 329 39081
rect 71 38978 82 39070
rect 318 38978 329 39070
rect 71 38967 329 38978
rect 71 38921 174 38967
rect 220 38921 329 38967
rect 71 38910 329 38921
rect 71 38818 82 38910
rect 318 38818 329 38910
rect 71 38807 329 38818
rect 71 38761 174 38807
rect 220 38761 329 38807
rect 71 38750 329 38761
rect 71 38658 82 38750
rect 318 38658 329 38750
rect 71 38647 329 38658
rect 71 38601 174 38647
rect 220 38601 329 38647
rect 71 38590 329 38601
rect 71 38498 82 38590
rect 318 38498 329 38590
rect 71 38487 329 38498
rect 71 38441 174 38487
rect 220 38441 329 38487
rect 71 38430 329 38441
rect 71 38338 82 38430
rect 318 38338 329 38430
rect 71 38327 329 38338
rect 71 38281 174 38327
rect 220 38281 329 38327
rect 71 38270 329 38281
rect 71 38178 82 38270
rect 318 38178 329 38270
rect 71 38167 329 38178
rect 71 38121 174 38167
rect 220 38121 329 38167
rect 71 38110 329 38121
rect 71 38018 82 38110
rect 318 38018 329 38110
rect 71 38007 329 38018
rect 71 37961 174 38007
rect 220 37961 329 38007
rect 71 37950 329 37961
rect 71 37858 82 37950
rect 318 37858 329 37950
rect 71 37847 329 37858
rect 71 37801 174 37847
rect 220 37801 329 37847
rect 71 37790 329 37801
rect 71 37698 82 37790
rect 318 37698 329 37790
rect 71 37687 329 37698
rect 71 37641 174 37687
rect 220 37641 329 37687
rect 71 37630 329 37641
rect 71 37538 82 37630
rect 318 37538 329 37630
rect 71 37527 329 37538
rect 71 37481 174 37527
rect 220 37481 329 37527
rect 71 37470 329 37481
rect 71 37378 82 37470
rect 318 37378 329 37470
rect 71 37367 329 37378
rect 71 37321 174 37367
rect 220 37321 329 37367
rect 71 37310 329 37321
rect 71 37218 82 37310
rect 318 37218 329 37310
rect 71 37207 329 37218
rect 71 37161 174 37207
rect 220 37161 329 37207
rect 71 37150 329 37161
rect 71 37058 82 37150
rect 318 37058 329 37150
rect 71 37047 329 37058
rect 71 37001 174 37047
rect 220 37001 329 37047
rect 71 36990 329 37001
rect 71 36898 82 36990
rect 318 36898 329 36990
rect 71 36887 329 36898
rect 71 36841 174 36887
rect 220 36841 329 36887
rect 71 36830 329 36841
rect 71 36738 82 36830
rect 318 36738 329 36830
rect 71 36727 329 36738
rect 71 36681 174 36727
rect 220 36681 329 36727
rect 71 36670 329 36681
rect 71 36578 82 36670
rect 318 36578 329 36670
rect 71 36567 329 36578
rect 71 36521 174 36567
rect 220 36521 329 36567
rect 71 36510 329 36521
rect 71 36418 82 36510
rect 318 36418 329 36510
rect 71 36407 329 36418
rect 71 36361 174 36407
rect 220 36361 329 36407
rect 71 36350 329 36361
rect 71 36258 82 36350
rect 318 36258 329 36350
rect 71 36247 329 36258
rect 71 36201 174 36247
rect 220 36201 329 36247
rect 71 36190 329 36201
rect 71 36098 82 36190
rect 318 36098 329 36190
rect 71 36087 329 36098
rect 71 36041 174 36087
rect 220 36041 329 36087
rect 71 36030 329 36041
rect 71 35938 82 36030
rect 318 35938 329 36030
rect 71 35927 329 35938
rect 71 35881 174 35927
rect 220 35881 329 35927
rect 71 35870 329 35881
rect 71 35778 82 35870
rect 318 35778 329 35870
rect 71 35767 329 35778
rect 71 35721 174 35767
rect 220 35721 329 35767
rect 71 35710 329 35721
rect 71 35618 82 35710
rect 318 35618 329 35710
rect 71 35607 329 35618
rect 71 35561 174 35607
rect 220 35561 329 35607
rect 71 35550 329 35561
rect 71 35458 82 35550
rect 318 35458 329 35550
rect 71 35447 329 35458
rect 71 35401 174 35447
rect 220 35401 329 35447
rect 71 35390 329 35401
rect 71 35298 82 35390
rect 318 35298 329 35390
rect 71 35287 329 35298
rect 71 35241 174 35287
rect 220 35241 329 35287
rect 71 35230 329 35241
rect 71 35138 82 35230
rect 318 35138 329 35230
rect 71 35127 329 35138
rect 71 35081 174 35127
rect 220 35081 329 35127
rect 71 35070 329 35081
rect 71 34978 82 35070
rect 318 34978 329 35070
rect 71 34967 329 34978
rect 71 34921 174 34967
rect 220 34921 329 34967
rect 71 34910 329 34921
rect 71 34818 82 34910
rect 318 34818 329 34910
rect 71 34807 329 34818
rect 71 34761 174 34807
rect 220 34761 329 34807
rect 71 34750 329 34761
rect 71 34658 82 34750
rect 318 34658 329 34750
rect 71 34647 329 34658
rect 71 34601 174 34647
rect 220 34601 329 34647
rect 71 34590 329 34601
rect 71 34498 82 34590
rect 318 34498 329 34590
rect 71 34487 329 34498
rect 71 34441 174 34487
rect 220 34441 329 34487
rect 71 34430 329 34441
rect 71 34338 82 34430
rect 318 34338 329 34430
rect 71 34327 329 34338
rect 71 34281 174 34327
rect 220 34281 329 34327
rect 71 34270 329 34281
rect 71 34178 82 34270
rect 318 34178 329 34270
rect 71 34167 329 34178
rect 71 34121 174 34167
rect 220 34121 329 34167
rect 71 34110 329 34121
rect 71 34018 82 34110
rect 318 34018 329 34110
rect 71 34007 329 34018
rect 71 33961 174 34007
rect 220 33961 329 34007
rect 71 33950 329 33961
rect 71 33858 82 33950
rect 318 33858 329 33950
rect 71 33847 329 33858
rect 71 33801 174 33847
rect 220 33801 329 33847
rect 71 33790 329 33801
rect 71 33698 82 33790
rect 318 33698 329 33790
rect 71 33687 329 33698
rect 71 33641 174 33687
rect 220 33641 329 33687
rect 71 33630 329 33641
rect 71 33538 82 33630
rect 318 33538 329 33630
rect 71 33527 329 33538
rect 71 33481 174 33527
rect 220 33481 329 33527
rect 71 33470 329 33481
rect 71 33378 82 33470
rect 318 33378 329 33470
rect 71 33367 329 33378
rect 71 33321 174 33367
rect 220 33321 329 33367
rect 71 33310 329 33321
rect 71 33218 82 33310
rect 318 33218 329 33310
rect 71 33207 329 33218
rect 71 33161 174 33207
rect 220 33161 329 33207
rect 71 33150 329 33161
rect 71 33058 82 33150
rect 318 33058 329 33150
rect 71 33047 329 33058
rect 71 33001 174 33047
rect 220 33001 329 33047
rect 71 32990 329 33001
rect 71 32898 82 32990
rect 318 32898 329 32990
rect 71 32887 329 32898
rect 71 32841 174 32887
rect 220 32841 329 32887
rect 71 32830 329 32841
rect 71 32738 82 32830
rect 318 32738 329 32830
rect 71 32727 329 32738
rect 71 32681 174 32727
rect 220 32681 329 32727
rect 71 32670 329 32681
rect 71 32578 82 32670
rect 318 32578 329 32670
rect 71 32567 329 32578
rect 71 32521 174 32567
rect 220 32521 329 32567
rect 71 32510 329 32521
rect 71 32418 82 32510
rect 318 32418 329 32510
rect 71 32407 329 32418
rect 71 32361 174 32407
rect 220 32361 329 32407
rect 71 32350 329 32361
rect 71 32258 82 32350
rect 318 32258 329 32350
rect 71 32247 329 32258
rect 71 32201 174 32247
rect 220 32201 329 32247
rect 71 32190 329 32201
rect 71 32098 82 32190
rect 318 32098 329 32190
rect 71 32087 329 32098
rect 71 32041 174 32087
rect 220 32041 329 32087
rect 71 32030 329 32041
rect 71 31938 82 32030
rect 318 31938 329 32030
rect 71 31927 329 31938
rect 71 31881 174 31927
rect 220 31881 329 31927
rect 71 31870 329 31881
rect 71 31778 82 31870
rect 318 31778 329 31870
rect 71 31767 329 31778
rect 71 31721 174 31767
rect 220 31721 329 31767
rect 71 31710 329 31721
rect 71 31618 82 31710
rect 318 31618 329 31710
rect 71 31607 329 31618
rect 71 31561 174 31607
rect 220 31561 329 31607
rect 71 31550 329 31561
rect 71 31458 82 31550
rect 318 31458 329 31550
rect 71 31447 329 31458
rect 71 31401 174 31447
rect 220 31401 329 31447
rect 71 31390 329 31401
rect 71 31298 82 31390
rect 318 31298 329 31390
rect 71 31287 329 31298
rect 71 31241 174 31287
rect 220 31241 329 31287
rect 71 31230 329 31241
rect 71 31138 82 31230
rect 318 31138 329 31230
rect 71 31127 329 31138
rect 71 31081 174 31127
rect 220 31081 329 31127
rect 71 31070 329 31081
rect 71 30978 82 31070
rect 318 30978 329 31070
rect 71 30967 329 30978
rect 71 30921 174 30967
rect 220 30921 329 30967
rect 71 30910 329 30921
rect 71 30818 82 30910
rect 318 30818 329 30910
rect 71 30807 329 30818
rect 71 30761 174 30807
rect 220 30761 329 30807
rect 71 30750 329 30761
rect 71 30658 82 30750
rect 318 30658 329 30750
rect 71 30647 329 30658
rect 71 30601 174 30647
rect 220 30601 329 30647
rect 71 30590 329 30601
rect 71 30498 82 30590
rect 318 30498 329 30590
rect 71 30487 329 30498
rect 71 30441 174 30487
rect 220 30441 329 30487
rect 71 30430 329 30441
rect 71 30338 82 30430
rect 318 30338 329 30430
rect 71 30327 329 30338
rect 71 30281 174 30327
rect 220 30281 329 30327
rect 71 30270 329 30281
rect 71 30178 82 30270
rect 318 30178 329 30270
rect 71 30167 329 30178
rect 71 30121 174 30167
rect 220 30121 329 30167
rect 71 30110 329 30121
rect 71 30018 82 30110
rect 318 30018 329 30110
rect 71 30007 329 30018
rect 71 29961 174 30007
rect 220 29961 329 30007
rect 71 29950 329 29961
rect 71 29858 82 29950
rect 318 29858 329 29950
rect 71 29847 329 29858
rect 71 29801 174 29847
rect 220 29801 329 29847
rect 71 29790 329 29801
rect 71 29698 82 29790
rect 318 29698 329 29790
rect 71 29687 329 29698
rect 71 29641 174 29687
rect 220 29641 329 29687
rect 71 29630 329 29641
rect 71 29538 82 29630
rect 318 29538 329 29630
rect 71 29527 329 29538
rect 71 29481 174 29527
rect 220 29481 329 29527
rect 71 29470 329 29481
rect 71 29378 82 29470
rect 318 29378 329 29470
rect 71 29367 329 29378
rect 71 29321 174 29367
rect 220 29321 329 29367
rect 71 29310 329 29321
rect 71 29218 82 29310
rect 318 29218 329 29310
rect 71 29207 329 29218
rect 71 29161 174 29207
rect 220 29161 329 29207
rect 71 29150 329 29161
rect 71 29058 82 29150
rect 318 29058 329 29150
rect 71 29047 329 29058
rect 71 29001 174 29047
rect 220 29001 329 29047
rect 71 28990 329 29001
rect 71 28898 82 28990
rect 318 28898 329 28990
rect 71 28887 329 28898
rect 71 28841 174 28887
rect 220 28841 329 28887
rect 71 28830 329 28841
rect 71 28738 82 28830
rect 318 28738 329 28830
rect 71 28727 329 28738
rect 71 28681 174 28727
rect 220 28681 329 28727
rect 71 28670 329 28681
rect 71 28578 82 28670
rect 318 28578 329 28670
rect 71 28567 329 28578
rect 71 28521 174 28567
rect 220 28521 329 28567
rect 71 28510 329 28521
rect 71 28418 82 28510
rect 318 28418 329 28510
rect 71 28407 329 28418
rect 71 28361 174 28407
rect 220 28361 329 28407
rect 71 28350 329 28361
rect 71 28258 82 28350
rect 318 28258 329 28350
rect 71 28247 329 28258
rect 71 28201 174 28247
rect 220 28201 329 28247
rect 71 28190 329 28201
rect 71 28098 82 28190
rect 318 28098 329 28190
rect 71 28087 329 28098
rect 71 28041 174 28087
rect 220 28041 329 28087
rect 71 28030 329 28041
rect 71 27938 82 28030
rect 318 27938 329 28030
rect 71 27927 329 27938
rect 71 27881 174 27927
rect 220 27881 329 27927
rect 71 27870 329 27881
rect 71 27778 82 27870
rect 318 27778 329 27870
rect 71 27767 329 27778
rect 71 27721 174 27767
rect 220 27721 329 27767
rect 71 27710 329 27721
rect 71 27618 82 27710
rect 318 27618 329 27710
rect 71 27607 329 27618
rect 71 27561 174 27607
rect 220 27561 329 27607
rect 71 27550 329 27561
rect 71 27458 82 27550
rect 318 27458 329 27550
rect 71 27447 329 27458
rect 71 27401 174 27447
rect 220 27401 329 27447
rect 71 27390 329 27401
rect 71 27298 82 27390
rect 318 27298 329 27390
rect 71 27287 329 27298
rect 71 27241 174 27287
rect 220 27241 329 27287
rect 71 27230 329 27241
rect 71 27138 82 27230
rect 318 27138 329 27230
rect 71 27127 329 27138
rect 71 27081 174 27127
rect 220 27081 329 27127
rect 71 27070 329 27081
rect 71 26978 82 27070
rect 318 26978 329 27070
rect 71 26967 329 26978
rect 71 26921 174 26967
rect 220 26921 329 26967
rect 71 26910 329 26921
rect 71 26818 82 26910
rect 318 26818 329 26910
rect 71 26807 329 26818
rect 71 26761 174 26807
rect 220 26761 329 26807
rect 71 26750 329 26761
rect 71 26658 82 26750
rect 318 26658 329 26750
rect 71 26647 329 26658
rect 71 26601 174 26647
rect 220 26601 329 26647
rect 71 26590 329 26601
rect 71 26498 82 26590
rect 318 26498 329 26590
rect 71 26487 329 26498
rect 71 26441 174 26487
rect 220 26441 329 26487
rect 71 26430 329 26441
rect 71 26338 82 26430
rect 318 26338 329 26430
rect 71 26327 329 26338
rect 71 26281 174 26327
rect 220 26281 329 26327
rect 71 26270 329 26281
rect 71 26178 82 26270
rect 318 26178 329 26270
rect 71 26167 329 26178
rect 71 26121 174 26167
rect 220 26121 329 26167
rect 71 26110 329 26121
rect 71 26018 82 26110
rect 318 26018 329 26110
rect 71 26007 329 26018
rect 71 25961 174 26007
rect 220 25961 329 26007
rect 71 25950 329 25961
rect 71 25858 82 25950
rect 318 25858 329 25950
rect 71 25847 329 25858
rect 71 25801 174 25847
rect 220 25801 329 25847
rect 71 25790 329 25801
rect 71 25698 82 25790
rect 318 25698 329 25790
rect 71 25687 329 25698
rect 71 25641 174 25687
rect 220 25641 329 25687
rect 71 25630 329 25641
rect 71 25538 82 25630
rect 318 25538 329 25630
rect 71 25527 329 25538
rect 71 25481 174 25527
rect 220 25481 329 25527
rect 71 25470 329 25481
rect 71 25378 82 25470
rect 318 25378 329 25470
rect 71 25367 329 25378
rect 71 25321 174 25367
rect 220 25321 329 25367
rect 71 25310 329 25321
rect 71 25218 82 25310
rect 318 25218 329 25310
rect 71 25207 329 25218
rect 71 25161 174 25207
rect 220 25161 329 25207
rect 71 25150 329 25161
rect 71 25058 82 25150
rect 318 25058 329 25150
rect 71 25047 329 25058
rect 71 25001 174 25047
rect 220 25001 329 25047
rect 71 24990 329 25001
rect 71 24898 82 24990
rect 318 24898 329 24990
rect 71 24887 329 24898
rect 71 24841 174 24887
rect 220 24841 329 24887
rect 71 24830 329 24841
rect 71 24738 82 24830
rect 318 24738 329 24830
rect 71 24727 329 24738
rect 71 24681 174 24727
rect 220 24681 329 24727
rect 71 24670 329 24681
rect 71 24578 82 24670
rect 318 24578 329 24670
rect 71 24567 329 24578
rect 71 24521 174 24567
rect 220 24521 329 24567
rect 71 24510 329 24521
rect 71 24418 82 24510
rect 318 24418 329 24510
rect 71 24407 329 24418
rect 71 24361 174 24407
rect 220 24361 329 24407
rect 71 24350 329 24361
rect 71 24258 82 24350
rect 318 24258 329 24350
rect 71 24247 329 24258
rect 71 24201 174 24247
rect 220 24201 329 24247
rect 71 24190 329 24201
rect 71 24098 82 24190
rect 318 24098 329 24190
rect 71 24087 329 24098
rect 71 24041 174 24087
rect 220 24041 329 24087
rect 71 24030 329 24041
rect 71 23938 82 24030
rect 318 23938 329 24030
rect 71 23927 329 23938
rect 71 23881 174 23927
rect 220 23881 329 23927
rect 71 23870 329 23881
rect 71 23778 82 23870
rect 318 23778 329 23870
rect 71 23767 329 23778
rect 71 23721 174 23767
rect 220 23721 329 23767
rect 71 23710 329 23721
rect 71 23618 82 23710
rect 318 23618 329 23710
rect 71 23607 329 23618
rect 71 23561 174 23607
rect 220 23561 329 23607
rect 71 23550 329 23561
rect 71 23458 82 23550
rect 318 23458 329 23550
rect 71 23447 329 23458
rect 71 23401 174 23447
rect 220 23401 329 23447
rect 71 23390 329 23401
rect 71 23298 82 23390
rect 318 23298 329 23390
rect 71 23287 329 23298
rect 71 23241 174 23287
rect 220 23241 329 23287
rect 71 23230 329 23241
rect 71 23138 82 23230
rect 318 23138 329 23230
rect 71 23127 329 23138
rect 71 23081 174 23127
rect 220 23081 329 23127
rect 71 23070 329 23081
rect 71 22978 82 23070
rect 318 22978 329 23070
rect 71 22967 329 22978
rect 71 22921 174 22967
rect 220 22921 329 22967
rect 71 22910 329 22921
rect 71 22818 82 22910
rect 318 22818 329 22910
rect 71 22807 329 22818
rect 71 22761 174 22807
rect 220 22761 329 22807
rect 71 22750 329 22761
rect 71 22658 82 22750
rect 318 22658 329 22750
rect 71 22647 329 22658
rect 71 22601 174 22647
rect 220 22601 329 22647
rect 71 22590 329 22601
rect 71 22498 82 22590
rect 318 22498 329 22590
rect 71 22487 329 22498
rect 71 22441 174 22487
rect 220 22441 329 22487
rect 71 22430 329 22441
rect 71 22338 82 22430
rect 318 22338 329 22430
rect 71 22327 329 22338
rect 71 22281 174 22327
rect 220 22281 329 22327
rect 71 22270 329 22281
rect 71 22178 82 22270
rect 318 22178 329 22270
rect 71 22167 329 22178
rect 71 22121 174 22167
rect 220 22121 329 22167
rect 71 22110 329 22121
rect 71 22018 82 22110
rect 318 22018 329 22110
rect 71 22007 329 22018
rect 71 21961 174 22007
rect 220 21961 329 22007
rect 71 21950 329 21961
rect 71 21858 82 21950
rect 318 21858 329 21950
rect 71 21847 329 21858
rect 71 21801 174 21847
rect 220 21801 329 21847
rect 71 21790 329 21801
rect 71 21698 82 21790
rect 318 21698 329 21790
rect 71 21687 329 21698
rect 71 21641 174 21687
rect 220 21641 329 21687
rect 71 21630 329 21641
rect 71 21538 82 21630
rect 318 21538 329 21630
rect 71 21527 329 21538
rect 71 21481 174 21527
rect 220 21481 329 21527
rect 71 21470 329 21481
rect 71 21378 82 21470
rect 318 21378 329 21470
rect 71 21367 329 21378
rect 71 21321 174 21367
rect 220 21321 329 21367
rect 71 21310 329 21321
rect 71 21218 82 21310
rect 318 21218 329 21310
rect 71 21207 329 21218
rect 71 21161 174 21207
rect 220 21161 329 21207
rect 71 21150 329 21161
rect 71 21058 82 21150
rect 318 21058 329 21150
rect 71 21047 329 21058
rect 71 21001 174 21047
rect 220 21001 329 21047
rect 71 20990 329 21001
rect 71 20898 82 20990
rect 318 20898 329 20990
rect 71 20887 329 20898
rect 71 20841 174 20887
rect 220 20841 329 20887
rect 71 20830 329 20841
rect 71 20738 82 20830
rect 318 20738 329 20830
rect 71 20727 329 20738
rect 71 20681 174 20727
rect 220 20681 329 20727
rect 71 20670 329 20681
rect 71 20578 82 20670
rect 318 20578 329 20670
rect 71 20567 329 20578
rect 71 20521 174 20567
rect 220 20521 329 20567
rect 71 20510 329 20521
rect 71 20418 82 20510
rect 318 20418 329 20510
rect 71 20407 329 20418
rect 71 20361 174 20407
rect 220 20361 329 20407
rect 71 20350 329 20361
rect 71 20258 82 20350
rect 318 20258 329 20350
rect 71 20247 329 20258
rect 71 20201 174 20247
rect 220 20201 329 20247
rect 71 20190 329 20201
rect 71 20098 82 20190
rect 318 20098 329 20190
rect 71 20087 329 20098
rect 71 20041 174 20087
rect 220 20041 329 20087
rect 71 20030 329 20041
rect 71 19938 82 20030
rect 318 19938 329 20030
rect 71 19927 329 19938
rect 71 19881 174 19927
rect 220 19881 329 19927
rect 71 19870 329 19881
rect 71 19778 82 19870
rect 318 19778 329 19870
rect 71 19767 329 19778
rect 71 19721 174 19767
rect 220 19721 329 19767
rect 71 19710 329 19721
rect 71 19618 82 19710
rect 318 19618 329 19710
rect 71 19607 329 19618
rect 71 19561 174 19607
rect 220 19561 329 19607
rect 71 19550 329 19561
rect 71 19458 82 19550
rect 318 19458 329 19550
rect 71 19447 329 19458
rect 71 19401 174 19447
rect 220 19401 329 19447
rect 71 19390 329 19401
rect 71 19298 82 19390
rect 318 19298 329 19390
rect 71 19287 329 19298
rect 71 19241 174 19287
rect 220 19241 329 19287
rect 71 19230 329 19241
rect 71 19138 82 19230
rect 318 19138 329 19230
rect 71 19127 329 19138
rect 71 19081 174 19127
rect 220 19081 329 19127
rect 71 19070 329 19081
rect 71 18978 82 19070
rect 318 18978 329 19070
rect 71 18967 329 18978
rect 71 18921 174 18967
rect 220 18921 329 18967
rect 71 18910 329 18921
rect 71 18818 82 18910
rect 318 18818 329 18910
rect 71 18807 329 18818
rect 71 18761 174 18807
rect 220 18761 329 18807
rect 71 18750 329 18761
rect 71 18658 82 18750
rect 318 18658 329 18750
rect 71 18647 329 18658
rect 71 18601 174 18647
rect 220 18601 329 18647
rect 71 18590 329 18601
rect 71 18498 82 18590
rect 318 18498 329 18590
rect 71 18487 329 18498
rect 71 18441 174 18487
rect 220 18441 329 18487
rect 71 18430 329 18441
rect 71 18338 82 18430
rect 318 18338 329 18430
rect 71 18327 329 18338
rect 71 18281 174 18327
rect 220 18281 329 18327
rect 71 18270 329 18281
rect 71 18178 82 18270
rect 318 18178 329 18270
rect 71 18167 329 18178
rect 71 18121 174 18167
rect 220 18121 329 18167
rect 71 18110 329 18121
rect 71 18018 82 18110
rect 318 18018 329 18110
rect 71 18007 329 18018
rect 71 17961 174 18007
rect 220 17961 329 18007
rect 71 17950 329 17961
rect 71 17858 82 17950
rect 318 17858 329 17950
rect 71 17847 329 17858
rect 71 17801 174 17847
rect 220 17801 329 17847
rect 71 17790 329 17801
rect 71 17698 82 17790
rect 318 17698 329 17790
rect 71 17687 329 17698
rect 71 17641 174 17687
rect 220 17641 329 17687
rect 71 17630 329 17641
rect 71 17538 82 17630
rect 318 17538 329 17630
rect 71 17527 329 17538
rect 71 17481 174 17527
rect 220 17481 329 17527
rect 71 17470 329 17481
rect 71 17378 82 17470
rect 318 17378 329 17470
rect 71 17367 329 17378
rect 71 17321 174 17367
rect 220 17321 329 17367
rect 71 17310 329 17321
rect 71 17218 82 17310
rect 318 17218 329 17310
rect 71 17207 329 17218
rect 71 17161 174 17207
rect 220 17161 329 17207
rect 71 17150 329 17161
rect 71 17058 82 17150
rect 318 17058 329 17150
rect 71 17047 329 17058
rect 71 17001 174 17047
rect 220 17001 329 17047
rect 71 16990 329 17001
rect 71 16898 82 16990
rect 318 16898 329 16990
rect 71 16887 329 16898
rect 71 16841 174 16887
rect 220 16841 329 16887
rect 71 16830 329 16841
rect 71 16738 82 16830
rect 318 16738 329 16830
rect 71 16727 329 16738
rect 71 16681 174 16727
rect 220 16681 329 16727
rect 71 16670 329 16681
rect 71 16578 82 16670
rect 318 16578 329 16670
rect 71 16567 329 16578
rect 71 16521 174 16567
rect 220 16521 329 16567
rect 71 16510 329 16521
rect 71 16418 82 16510
rect 318 16418 329 16510
rect 71 16407 329 16418
rect 71 16361 174 16407
rect 220 16361 329 16407
rect 71 16350 329 16361
rect 71 16258 82 16350
rect 318 16258 329 16350
rect 71 16247 329 16258
rect 71 16201 174 16247
rect 220 16201 329 16247
rect 71 16190 329 16201
rect 71 16098 82 16190
rect 318 16098 329 16190
rect 71 16087 329 16098
rect 71 16041 174 16087
rect 220 16041 329 16087
rect 71 16030 329 16041
rect 71 15938 82 16030
rect 318 15938 329 16030
rect 71 15927 329 15938
rect 71 15881 174 15927
rect 220 15881 329 15927
rect 71 15870 329 15881
rect 71 15778 82 15870
rect 318 15778 329 15870
rect 71 15767 329 15778
rect 71 15721 174 15767
rect 220 15721 329 15767
rect 71 15710 329 15721
rect 71 15618 82 15710
rect 318 15618 329 15710
rect 71 15607 329 15618
rect 71 15561 174 15607
rect 220 15561 329 15607
rect 71 15550 329 15561
rect 71 15458 82 15550
rect 318 15458 329 15550
rect 71 15447 329 15458
rect 71 15401 174 15447
rect 220 15401 329 15447
rect 71 15390 329 15401
rect 71 15298 82 15390
rect 318 15298 329 15390
rect 71 15287 329 15298
rect 71 15241 174 15287
rect 220 15241 329 15287
rect 71 15230 329 15241
rect 71 15138 82 15230
rect 318 15138 329 15230
rect 71 15127 329 15138
rect 71 15081 174 15127
rect 220 15081 329 15127
rect 71 15070 329 15081
rect 71 14978 82 15070
rect 318 14978 329 15070
rect 71 14967 329 14978
rect 71 14921 174 14967
rect 220 14921 329 14967
rect 71 14910 329 14921
rect 71 14818 82 14910
rect 318 14818 329 14910
rect 71 14807 329 14818
rect 71 14761 174 14807
rect 220 14761 329 14807
rect 71 14750 329 14761
rect 71 14658 82 14750
rect 318 14658 329 14750
rect 71 14647 329 14658
rect 71 14601 174 14647
rect 220 14601 329 14647
rect 71 14590 329 14601
rect 71 14498 82 14590
rect 318 14498 329 14590
rect 71 14487 329 14498
rect 71 14441 174 14487
rect 220 14441 329 14487
rect 71 14430 329 14441
rect 71 14338 82 14430
rect 318 14338 329 14430
rect 71 14327 329 14338
rect 71 14281 174 14327
rect 220 14281 329 14327
rect 71 14270 329 14281
rect 71 14178 82 14270
rect 318 14178 329 14270
rect 71 14167 329 14178
rect 71 14121 174 14167
rect 220 14121 329 14167
rect 71 14110 329 14121
rect 71 14018 82 14110
rect 318 14018 329 14110
rect 71 14007 329 14018
rect 71 13961 174 14007
rect 220 13961 329 14007
rect 71 13950 329 13961
rect 71 13858 82 13950
rect 318 13858 329 13950
rect 71 13847 329 13858
rect 71 13801 174 13847
rect 220 13801 329 13847
rect 71 13790 329 13801
rect 71 13698 82 13790
rect 318 13698 329 13790
rect 71 13687 329 13698
rect 71 13641 174 13687
rect 220 13641 329 13687
rect 71 13630 329 13641
rect 71 13538 82 13630
rect 318 13538 329 13630
rect 71 13527 329 13538
rect 71 13481 174 13527
rect 220 13481 329 13527
rect 71 13470 329 13481
rect 71 13356 82 13470
rect -32 13276 82 13356
rect 318 13356 329 13470
rect 375 13356 432 69708
rect 318 13276 432 13356
rect -32 13262 432 13276
rect -32 13231 130 13262
rect -32 13185 25 13231
rect 71 13185 130 13231
rect -32 13122 130 13185
rect 270 13231 432 13262
rect 270 13185 329 13231
rect 375 13185 432 13231
rect 270 13122 432 13185
rect -32 13108 432 13122
<< via1 >>
rect 130 64890 286 64942
rect 130 64778 286 64830
rect 130 64681 174 64718
rect 174 64681 220 64718
rect 220 64681 286 64718
rect 130 64666 286 64681
rect 130 64567 286 64606
rect 130 64554 174 64567
rect 174 64554 220 64567
rect 220 64554 286 64567
rect 130 64442 286 64494
rect 130 64361 174 64382
rect 174 64361 220 64382
rect 220 64361 286 64382
rect 130 64330 286 64361
rect 130 64247 286 64270
rect 130 64218 174 64247
rect 174 64218 220 64247
rect 220 64218 286 64247
rect 130 64106 286 64158
rect 130 64041 174 64046
rect 174 64041 220 64046
rect 220 64041 286 64046
rect 130 63994 286 64041
rect 130 63927 286 63934
rect 130 63882 174 63927
rect 174 63882 220 63927
rect 220 63882 286 63927
rect 130 63770 286 63822
rect 130 63658 286 63710
rect 127 50487 179 50536
rect 127 50484 174 50487
rect 174 50484 179 50487
rect 239 50484 291 50536
rect 127 50372 179 50424
rect 239 50372 291 50424
rect 127 50281 174 50312
rect 174 50281 179 50312
rect 127 50260 179 50281
rect 239 50260 291 50312
rect 127 50167 179 50200
rect 127 50148 174 50167
rect 174 50148 179 50167
rect 239 50148 291 50200
rect 127 50036 179 50088
rect 239 50036 291 50088
rect 127 49961 174 49976
rect 174 49961 179 49976
rect 127 49924 179 49961
rect 239 49924 291 49976
rect 127 49847 179 49864
rect 127 49812 174 49847
rect 174 49812 179 49847
rect 239 49812 291 49864
rect 127 49700 179 49752
rect 239 49700 291 49752
rect 127 49588 179 49640
rect 239 49588 291 49640
rect 127 49527 179 49528
rect 127 49481 174 49527
rect 174 49481 179 49527
rect 127 49476 179 49481
rect 239 49476 291 49528
rect 127 49367 179 49416
rect 127 49364 174 49367
rect 174 49364 179 49367
rect 239 49364 291 49416
rect 127 49252 179 49304
rect 239 49252 291 49304
<< metal2 >>
rect 118 65000 298 69769
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 118 50600 298 63600
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
rect 118 13275 298 49200
<< via2 >>
rect 128 64942 288 64944
rect 128 64890 130 64942
rect 130 64890 286 64942
rect 286 64890 288 64942
rect 128 64888 288 64890
rect 128 64830 288 64832
rect 128 64778 130 64830
rect 130 64778 286 64830
rect 286 64778 288 64830
rect 128 64776 288 64778
rect 128 64718 288 64720
rect 128 64666 130 64718
rect 130 64666 286 64718
rect 286 64666 288 64718
rect 128 64664 288 64666
rect 128 64606 288 64608
rect 128 64554 130 64606
rect 130 64554 286 64606
rect 286 64554 288 64606
rect 128 64552 288 64554
rect 128 64494 288 64496
rect 128 64442 130 64494
rect 130 64442 286 64494
rect 286 64442 288 64494
rect 128 64440 288 64442
rect 128 64382 288 64384
rect 128 64330 130 64382
rect 130 64330 286 64382
rect 286 64330 288 64382
rect 128 64328 288 64330
rect 128 64270 288 64272
rect 128 64218 130 64270
rect 130 64218 286 64270
rect 286 64218 288 64270
rect 128 64216 288 64218
rect 128 64158 288 64160
rect 128 64106 130 64158
rect 130 64106 286 64158
rect 286 64106 288 64158
rect 128 64104 288 64106
rect 128 64046 288 64048
rect 128 63994 130 64046
rect 130 63994 286 64046
rect 286 63994 288 64046
rect 128 63992 288 63994
rect 128 63934 288 63936
rect 128 63882 130 63934
rect 130 63882 286 63934
rect 286 63882 288 63934
rect 128 63880 288 63882
rect 128 63822 288 63824
rect 128 63770 130 63822
rect 130 63770 286 63822
rect 286 63770 288 63822
rect 128 63768 288 63770
rect 128 63710 288 63712
rect 128 63658 130 63710
rect 130 63658 286 63710
rect 286 63658 288 63710
rect 128 63656 288 63658
rect 125 50536 181 50538
rect 125 50484 127 50536
rect 127 50484 179 50536
rect 179 50484 181 50536
rect 125 50482 181 50484
rect 237 50536 293 50538
rect 237 50484 239 50536
rect 239 50484 291 50536
rect 291 50484 293 50536
rect 237 50482 293 50484
rect 125 50424 181 50426
rect 125 50372 127 50424
rect 127 50372 179 50424
rect 179 50372 181 50424
rect 125 50370 181 50372
rect 237 50424 293 50426
rect 237 50372 239 50424
rect 239 50372 291 50424
rect 291 50372 293 50424
rect 237 50370 293 50372
rect 125 50312 181 50314
rect 125 50260 127 50312
rect 127 50260 179 50312
rect 179 50260 181 50312
rect 125 50258 181 50260
rect 237 50312 293 50314
rect 237 50260 239 50312
rect 239 50260 291 50312
rect 291 50260 293 50312
rect 237 50258 293 50260
rect 125 50200 181 50202
rect 125 50148 127 50200
rect 127 50148 179 50200
rect 179 50148 181 50200
rect 125 50146 181 50148
rect 237 50200 293 50202
rect 237 50148 239 50200
rect 239 50148 291 50200
rect 291 50148 293 50200
rect 237 50146 293 50148
rect 125 50088 181 50090
rect 125 50036 127 50088
rect 127 50036 179 50088
rect 179 50036 181 50088
rect 125 50034 181 50036
rect 237 50088 293 50090
rect 237 50036 239 50088
rect 239 50036 291 50088
rect 291 50036 293 50088
rect 237 50034 293 50036
rect 125 49976 181 49978
rect 125 49924 127 49976
rect 127 49924 179 49976
rect 179 49924 181 49976
rect 125 49922 181 49924
rect 237 49976 293 49978
rect 237 49924 239 49976
rect 239 49924 291 49976
rect 291 49924 293 49976
rect 237 49922 293 49924
rect 125 49864 181 49866
rect 125 49812 127 49864
rect 127 49812 179 49864
rect 179 49812 181 49864
rect 125 49810 181 49812
rect 237 49864 293 49866
rect 237 49812 239 49864
rect 239 49812 291 49864
rect 291 49812 293 49864
rect 237 49810 293 49812
rect 125 49752 181 49754
rect 125 49700 127 49752
rect 127 49700 179 49752
rect 179 49700 181 49752
rect 125 49698 181 49700
rect 237 49752 293 49754
rect 237 49700 239 49752
rect 239 49700 291 49752
rect 291 49700 293 49752
rect 237 49698 293 49700
rect 125 49640 181 49642
rect 125 49588 127 49640
rect 127 49588 179 49640
rect 179 49588 181 49640
rect 125 49586 181 49588
rect 237 49640 293 49642
rect 237 49588 239 49640
rect 239 49588 291 49640
rect 291 49588 293 49640
rect 237 49586 293 49588
rect 125 49528 181 49530
rect 125 49476 127 49528
rect 127 49476 179 49528
rect 179 49476 181 49528
rect 125 49474 181 49476
rect 237 49528 293 49530
rect 237 49476 239 49528
rect 239 49476 291 49528
rect 291 49476 293 49528
rect 237 49474 293 49476
rect 125 49416 181 49418
rect 125 49364 127 49416
rect 127 49364 179 49416
rect 179 49364 181 49416
rect 125 49362 181 49364
rect 237 49416 293 49418
rect 237 49364 239 49416
rect 239 49364 291 49416
rect 291 49364 293 49416
rect 237 49362 293 49364
rect 125 49304 181 49306
rect 125 49252 127 49304
rect 127 49252 179 49304
rect 179 49252 181 49304
rect 125 49250 181 49252
rect 237 49304 293 49306
rect 237 49252 239 49304
rect 239 49252 291 49304
rect 291 49252 293 49304
rect 237 49250 293 49252
<< metal3 >>
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
use POLY_FILL  POLY_FILL_0
array 0 0 0 0 351 160
timestamp 1764353313
transform 1 0 82 0 1 13462
box 0 0 1 1
<< labels >>
rlabel metal3 s 208 50023 208 50023 4 VSS
port 1 nsew
rlabel metal3 s 207 64258 207 64258 4 VSS
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 400 70000
string GDS_END 14026650
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 13941104
<< end >>
