magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< pwell >>
rect 597 223 1973 3135
<< mvndiff >>
rect 597 3069 685 3135
rect 597 1801 610 3069
rect 656 1801 685 3069
rect 597 1735 685 1801
rect 1885 3069 1973 3135
rect 1885 1801 1914 3069
rect 1960 1801 1973 3069
rect 1885 1735 1973 1801
rect 597 1557 685 1623
rect 597 289 610 1557
rect 656 289 685 1557
rect 597 223 685 289
rect 1885 1557 1973 1623
rect 1885 289 1914 1557
rect 1960 289 1973 1557
rect 1885 223 1973 289
<< mvndiffc >>
rect 610 1801 656 3069
rect 1914 1801 1960 3069
rect 610 289 656 1557
rect 1914 289 1960 1557
<< mvnmoscap >>
rect 685 1735 1885 3135
rect 685 223 1885 1623
<< polysilicon >>
rect 685 3214 1885 3227
rect 685 3168 745 3214
rect 1825 3168 1885 3214
rect 685 3135 1885 3168
rect 685 1702 1885 1735
rect 685 1656 745 1702
rect 1825 1656 1885 1702
rect 685 1623 1885 1656
rect 685 190 1885 223
rect 685 144 745 190
rect 1825 144 1885 190
rect 685 131 1885 144
<< polycontact >>
rect 745 3168 1825 3214
rect 745 1656 1825 1702
rect 745 144 1825 190
<< metal1 >>
rect 310 3285 2260 3485
rect 310 3069 667 3285
rect 727 3214 1843 3225
rect 727 3168 745 3214
rect 1825 3168 1843 3214
rect 727 3161 1088 3168
rect 1140 3161 1220 3168
rect 1272 3161 1352 3168
rect 1404 3161 1843 3168
rect 727 3157 1843 3161
rect 310 1801 610 3069
rect 656 1801 667 3069
rect 310 1557 667 1801
rect 785 1713 1785 3157
rect 1903 3069 2260 3285
rect 1903 1801 1914 3069
rect 1960 1801 2260 3069
rect 727 1702 1843 1713
rect 727 1656 745 1702
rect 1825 1656 1843 1702
rect 727 1645 1843 1656
rect 310 289 610 1557
rect 656 289 667 1557
rect 310 73 667 289
rect 785 201 1785 1645
rect 1903 1557 2260 1801
rect 1903 289 1914 1557
rect 1960 289 2260 1557
rect 727 197 1843 201
rect 727 190 1088 197
rect 1140 190 1220 197
rect 1272 190 1352 197
rect 1404 190 1843 197
rect 727 144 745 190
rect 1825 144 1843 190
rect 727 133 1843 144
rect 1903 73 2260 289
rect 310 -127 2260 73
<< via1 >>
rect 1088 3168 1140 3213
rect 1220 3168 1272 3213
rect 1352 3168 1404 3213
rect 1088 3161 1140 3168
rect 1220 3161 1272 3168
rect 1352 3161 1404 3168
rect 1088 190 1140 197
rect 1220 190 1272 197
rect 1352 190 1404 197
rect 1088 145 1140 190
rect 1220 145 1272 190
rect 1352 145 1404 190
<< metal2 >>
rect 1076 3213 1427 3485
rect 1076 3161 1088 3213
rect 1140 3161 1220 3213
rect 1272 3161 1352 3213
rect 1404 3161 1427 3213
rect 1076 197 1427 3161
rect 1076 145 1088 197
rect 1140 145 1220 197
rect 1272 145 1352 197
rect 1404 145 1427 197
rect 1076 -127 1427 145
<< properties >>
string GDS_END 54010690
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 54003006
<< end >>
