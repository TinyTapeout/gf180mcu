magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect -1789 9497 11222 10481
rect -1789 -266 -560 9497
rect 10028 -266 11222 9497
rect -1789 -834 11222 -266
<< psubdiff >>
rect -528 8756 9996 9430
rect -528 8372 9406 8756
rect -528 -174 -486 8372
rect -140 8195 9406 8372
rect 9586 8372 9996 8756
rect -140 -35 -118 8195
rect 9586 -35 9608 8372
rect -140 -57 9608 -35
rect -140 -174 208 -57
rect -528 -197 208 -174
rect 9278 -174 9608 -57
rect 9954 -174 9996 8372
rect 9278 -197 9996 -174
rect -528 -219 9996 -197
<< nsubdiff >>
rect -1707 10362 11139 10398
rect -1707 9616 -421 10362
rect 9925 9616 11139 10362
rect -1707 9580 11139 9616
rect -1707 8368 -643 9580
rect -1707 22 -1629 8368
rect -683 22 -643 8368
rect -1707 -83 -643 22
rect -1707 -729 -1629 -83
rect -683 -349 -643 -83
rect 10111 8368 11139 9580
rect 10111 22 10151 8368
rect 11097 22 11139 8368
rect 10111 -83 11139 22
rect 10111 -349 10151 -83
rect -683 -377 10151 -349
rect -683 -723 -413 -377
rect 9933 -723 10151 -377
rect -683 -729 10151 -723
rect 11097 -729 11139 -83
rect -1707 -751 11139 -729
<< psubdiffcont >>
rect -486 -174 -140 8372
rect 208 -197 9278 -57
rect 9608 -174 9954 8372
<< nsubdiffcont >>
rect -421 9616 9925 10362
rect -1629 22 -683 8368
rect -1629 -729 -683 -83
rect 10151 22 11097 8368
rect -413 -723 9933 -377
rect 10151 -729 11097 -83
<< metal1 >>
rect -432 10362 9936 10387
rect -432 9616 -421 10362
rect 9925 9616 9936 10362
rect -432 9591 9936 9616
rect -1658 8368 -654 8388
rect -1658 22 -1629 8368
rect -683 22 -654 8368
rect -1658 -83 -654 22
rect -1658 -729 -1629 -83
rect -683 -360 -654 -83
rect -517 8372 51 8396
rect -517 -174 -486 8372
rect -140 -46 51 8372
rect 9597 8372 9985 8383
rect 9597 -46 9608 8372
rect -140 -57 9608 -46
rect -140 -174 208 -57
rect -517 -197 208 -174
rect 9278 -174 9608 -57
rect 9954 -174 9985 8372
rect 9278 -197 9985 -174
rect -517 -208 9985 -197
rect 10122 8368 11126 8410
rect 10122 22 10151 8368
rect 11097 22 11126 8368
rect 10122 -83 11126 22
rect 10122 -360 10151 -83
rect -683 -377 10151 -360
rect -683 -723 -413 -377
rect 9933 -723 10151 -377
rect -683 -729 10151 -723
rect 11097 -729 11126 -83
rect -1658 -740 11126 -729
<< properties >>
string GDS_END 11077898
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 10823238
<< end >>
