magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect -1730 9497 11766 10481
rect -1730 -15 -500 9497
rect 10573 -15 11766 9497
rect -1730 -583 11766 -15
<< psubdiff >>
rect -458 8756 10536 9430
rect -458 8289 -118 8756
rect -458 65 -390 8289
rect -156 322 -118 8289
rect 10146 8322 10536 8756
rect 10146 8300 10541 8322
rect 10146 322 10173 8300
rect -156 294 10173 322
rect -156 65 29 294
rect -458 60 29 65
rect 10039 60 10173 294
rect -458 54 10173 60
rect 10519 54 10541 8300
rect -458 32 10541 54
<< nsubdiff >>
rect -1647 10362 11683 10398
rect -1647 9616 -436 10362
rect 10510 9616 11683 10362
rect -1647 9580 11683 9616
rect -1647 8368 -583 9580
rect -1647 -478 -1569 8368
rect -623 -98 -583 8368
rect 10656 8368 11683 9580
rect 10656 -98 10696 8368
rect -623 -126 10696 -98
rect -623 -472 -436 -126
rect 10510 -472 10696 -126
rect -623 -478 10696 -472
rect 11642 -478 11683 8368
rect -1647 -500 11683 -478
<< psubdiffcont >>
rect -390 65 -156 8289
rect 29 60 10039 294
rect 10173 54 10519 8300
<< nsubdiffcont >>
rect -436 9616 10510 10362
rect -1569 -478 -623 8368
rect -436 -472 10510 -126
rect 10696 -478 11642 8368
<< metal1 >>
rect -447 10362 10521 10387
rect -447 9616 -436 10362
rect 10510 9616 10521 10362
rect -447 9591 10521 9616
rect -1598 8368 -594 8388
rect -1598 -478 -1569 8368
rect -623 -109 -594 8368
rect -457 8289 111 8396
rect -457 65 -390 8289
rect -156 311 111 8289
rect 9962 8300 10530 8397
rect 9962 311 10173 8300
rect -156 294 10173 311
rect -156 65 29 294
rect -457 60 29 65
rect 10039 60 10173 294
rect -457 54 10173 60
rect 10519 54 10530 8300
rect -457 43 10530 54
rect 10666 8368 11670 8410
rect 10666 -109 10696 8368
rect -623 -126 10696 -109
rect -623 -472 -436 -126
rect 10510 -472 10696 -126
rect -623 -478 10696 -472
rect 11642 -478 11670 8368
rect -1598 -489 11670 -478
<< properties >>
string GDS_END 12530082
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 12271134
<< end >>
