magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect 0 12 1196 8252
<< mvpmos >>
rect 278 132 418 8132
<< mvpdiff >>
rect 120 8103 222 8132
rect 120 161 133 8103
rect 179 161 222 8103
rect 120 132 222 161
rect 974 8103 1076 8132
rect 974 161 1017 8103
rect 1063 161 1076 8103
rect 974 132 1076 161
<< mvpdiffc >>
rect 133 161 179 8103
rect 1017 161 1063 8103
<< polysilicon >>
rect 278 8132 418 8220
rect 278 44 418 132
<< mvpdiffres >>
rect 222 132 278 8132
rect 418 132 974 8132
<< metal1 >>
rect 133 8103 179 8132
rect 133 132 179 161
rect 1017 8103 1063 8132
rect 1017 132 1063 161
<< properties >>
string GDS_END 12687484
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 12675576
<< end >>
