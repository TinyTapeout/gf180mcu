magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect 15280 46078 15875 46628
<< nmos >>
rect 15581 45872 15637 45992
<< pmos >>
rect 15581 46164 15637 46404
<< ndiff >>
rect 15492 45956 15581 45992
rect 15492 45910 15506 45956
rect 15552 45910 15581 45956
rect 15492 45872 15581 45910
rect 15637 45955 15725 45992
rect 15637 45909 15666 45955
rect 15712 45909 15725 45955
rect 15637 45872 15725 45909
<< pdiff >>
rect 15493 46353 15581 46404
rect 15493 46213 15506 46353
rect 15552 46213 15581 46353
rect 15493 46164 15581 46213
rect 15637 46353 15725 46404
rect 15637 46213 15666 46353
rect 15712 46213 15725 46353
rect 15637 46164 15725 46213
<< ndiffc >>
rect 15506 45910 15552 45956
rect 15666 45909 15712 45955
<< pdiffc >>
rect 15506 46213 15552 46353
rect 15666 46213 15712 46353
<< psubdiff >>
rect 15366 45791 15789 45806
rect 15366 45745 15379 45791
rect 15425 45745 15730 45791
rect 15776 45745 15789 45791
rect 15366 45730 15789 45745
<< nsubdiff >>
rect 15366 46531 15789 46546
rect 15366 46485 15379 46531
rect 15425 46485 15730 46531
rect 15776 46485 15789 46531
rect 15366 46470 15789 46485
<< psubdiffcont >>
rect 15379 45745 15425 45791
rect 15730 45745 15776 45791
<< nsubdiffcont >>
rect 15379 46485 15425 46531
rect 15730 46485 15776 46531
<< polysilicon >>
rect 15581 46404 15637 46450
rect 15396 46204 15468 46254
rect 15396 46158 15409 46204
rect 15455 46158 15468 46204
rect 15396 46144 15468 46158
rect 15581 46144 15637 46164
rect 15396 46108 15637 46144
rect 15397 46022 15637 46058
rect 15397 46008 15469 46022
rect 15397 45962 15410 46008
rect 15456 45962 15469 46008
rect 15581 45992 15637 46022
rect 15397 45912 15469 45962
rect 15581 45828 15637 45872
<< polycontact >>
rect 15409 46158 15455 46204
rect 15410 45962 15456 46008
<< metal1 >>
rect 15366 46531 15789 46542
rect 15366 46485 15379 46531
rect 15425 46485 15730 46531
rect 15776 46485 15789 46531
rect 15366 46467 15789 46485
rect 15506 46353 15552 46401
rect 15409 46204 15455 46252
rect 15409 46110 15455 46158
rect 15410 46008 15456 46056
rect 15410 45914 15456 45962
rect 15506 45956 15552 46213
rect 15506 45876 15552 45910
rect 15666 46353 15712 46401
rect 15666 45955 15712 46213
rect 15666 45875 15712 45909
rect 15366 45791 15789 45810
rect 15366 45745 15379 45791
rect 15425 45745 15730 45791
rect 15776 45745 15789 45791
rect 15366 45734 15789 45745
<< properties >>
string GDS_END 10542116
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 10539680
<< end >>
