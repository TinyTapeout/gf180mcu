magic
tech gf180mcuD
timestamp 1764353313
<< properties >>
string GDS_END 13941060
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 13940864
<< end >>
