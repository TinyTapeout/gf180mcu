magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect 758 14151 14242 68951
<< obsm1 >>
rect -32 13108 15032 69957
<< metal2 >>
rect 3068 26874 3576 70000
rect 4204 26874 4712 70000
rect 5340 26874 5848 70000
rect 6476 26874 6984 70000
rect 8016 26874 8524 70000
rect 9152 26874 9660 70000
rect 10288 26874 10796 70000
rect 11424 26874 11932 70000
<< obsm2 >>
rect 0 26814 3008 69678
rect 3636 26814 4144 69678
rect 4772 26814 5280 69678
rect 5908 26814 6416 69678
rect 7044 26814 7956 69678
rect 8584 26814 9092 69678
rect 9720 26814 10228 69678
rect 10856 26814 11364 69678
rect 11992 26814 15000 69678
rect 0 0 15000 26814
<< obsm3 >>
rect 0 0 15000 69678
<< obsm4 >>
rect 0 0 15000 69678
<< metal5 >>
rect 0 68400 1000 69678
rect 0 66800 1000 68200
rect 0 65200 1000 66600
rect 0 63600 1000 65000
rect 0 62000 1000 63400
rect 0 60400 1000 61800
rect 0 58800 1000 60200
rect 0 57200 1000 58600
rect 0 55600 1000 57000
rect 0 54000 1000 55400
rect 0 52400 1000 53800
rect 0 50800 1000 52200
rect 0 49200 1000 50600
rect 0 46000 1000 49000
rect 0 42800 1000 45800
rect 0 41200 1000 42600
rect 0 39600 1000 41000
rect 0 36400 1000 39400
rect 0 33200 1000 36200
rect 0 30000 1000 33000
rect 0 26800 1000 29800
rect 0 25200 1000 26600
rect 0 23600 1000 25000
rect 0 20400 1000 23400
rect 0 17200 1000 20200
rect 0 14000 1000 17000
rect 14000 68400 15000 69678
rect 14000 66800 15000 68200
rect 14000 65200 15000 66600
rect 14000 63600 15000 65000
rect 14000 62000 15000 63400
rect 14000 60400 15000 61800
rect 14000 58800 15000 60200
rect 14000 57200 15000 58600
rect 14000 55600 15000 57000
rect 14000 54000 15000 55400
rect 14000 52400 15000 53800
rect 14000 50800 15000 52200
rect 14000 49200 15000 50600
rect 14000 46000 15000 49000
rect 14000 42800 15000 45800
rect 14000 41200 15000 42600
rect 14000 39600 15000 41000
rect 14000 36400 15000 39400
rect 14000 33200 15000 36200
rect 14000 30000 15000 33000
rect 14000 26800 15000 29800
rect 14000 25200 15000 26600
rect 14000 23600 15000 25000
rect 14000 20400 15000 23400
rect 14000 17200 15000 20200
rect 14000 14000 15000 17000
rect 1500 400 13500 12400
<< obsm5 >>
rect 1120 13880 13880 69678
rect 700 12520 14300 13880
rect 700 280 1380 12520
rect 13620 280 14300 12520
rect 700 0 14300 280
<< labels >>
rlabel metal2 s 3068 26874 3576 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 4204 26874 4712 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 5340 26874 5848 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 6476 26874 6984 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 8016 26874 8524 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 9152 26874 9660 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 10288 26874 10796 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal2 s 11424 26874 11932 70000 6 ASIG5V
port 1 nsew signal bidirectional
rlabel metal5 s 0 66800 1000 68200 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 58800 1000 60200 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 55600 1000 57000 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 54000 1000 55400 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 52400 1000 53800 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 42800 1000 45800 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 41200 1000 42600 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 36400 1000 39400 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 33200 1000 36200 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 30000 1000 33000 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 26800 1000 29800 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 23600 1000 25000 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 66800 15000 68200 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 58800 15000 60200 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 55600 15000 57000 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 54000 15000 55400 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 52400 15000 53800 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 42800 15000 45800 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 41200 15000 42600 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 36400 15000 39400 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 33200 15000 36200 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 30000 15000 33000 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 26800 15000 29800 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 14000 23600 15000 25000 6 DVDD
port 2 nsew power bidirectional
rlabel metal5 s 0 17200 1000 20200 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 65200 1000 66600 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 68400 1000 69678 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 46000 1000 49000 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 57200 1000 58600 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 60400 1000 61800 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 39600 1000 41000 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 20400 1000 23400 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 25200 1000 26600 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 14000 1000 17000 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 17200 15000 20200 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 65200 15000 66600 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 68400 15000 69678 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 46000 15000 49000 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 57200 15000 58600 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 60400 15000 61800 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 39600 15000 41000 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 20400 15000 23400 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 25200 15000 26600 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 14000 14000 15000 17000 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 1500 400 13500 12400 6 DVSS
port 3 nsew ground bidirectional
rlabel metal5 s 0 62000 1000 63400 6 VDD
port 4 nsew power bidirectional
rlabel metal5 s 0 50800 1000 52200 6 VDD
port 4 nsew power bidirectional
rlabel metal5 s 14000 62000 15000 63400 6 VDD
port 4 nsew power bidirectional
rlabel metal5 s 14000 50800 15000 52200 6 VDD
port 4 nsew power bidirectional
rlabel metal5 s 0 63600 1000 65000 6 VSS
port 5 nsew ground bidirectional
rlabel metal5 s 0 49200 1000 50600 6 VSS
port 5 nsew ground bidirectional
rlabel metal5 s 14000 63600 15000 65000 6 VSS
port 5 nsew ground bidirectional
rlabel metal5 s 14000 49200 15000 50600 6 VSS
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string LEFclass PAD INOUT
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 10215176
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 10203210
<< end >>
