magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect -13 1870 695 2578
rect 1136 1870 1844 2578
rect -13 970 695 1678
rect 1136 970 1844 1678
<< nsubdiff >>
rect 73 2479 609 2492
rect 73 2433 86 2479
rect 132 2433 202 2479
rect 248 2433 318 2479
rect 364 2433 434 2479
rect 480 2433 550 2479
rect 596 2433 609 2479
rect 73 2420 609 2433
rect 73 2363 145 2420
rect 73 2317 86 2363
rect 132 2317 145 2363
rect 537 2363 609 2420
rect 73 2247 145 2317
rect 73 2201 86 2247
rect 132 2201 145 2247
rect 73 2131 145 2201
rect 73 2085 86 2131
rect 132 2085 145 2131
rect 537 2317 550 2363
rect 596 2317 609 2363
rect 537 2247 609 2317
rect 537 2201 550 2247
rect 596 2201 609 2247
rect 537 2131 609 2201
rect 73 2028 145 2085
rect 537 2085 550 2131
rect 596 2085 609 2131
rect 537 2028 609 2085
rect 73 2015 609 2028
rect 73 1969 86 2015
rect 132 1969 202 2015
rect 248 1969 318 2015
rect 364 1969 434 2015
rect 480 1969 550 2015
rect 596 1969 609 2015
rect 73 1956 609 1969
rect 1222 2479 1758 2492
rect 1222 2433 1235 2479
rect 1281 2433 1351 2479
rect 1397 2433 1467 2479
rect 1513 2433 1583 2479
rect 1629 2433 1699 2479
rect 1745 2433 1758 2479
rect 1222 2420 1758 2433
rect 1222 2363 1294 2420
rect 1222 2317 1235 2363
rect 1281 2317 1294 2363
rect 1686 2363 1758 2420
rect 1222 2247 1294 2317
rect 1222 2201 1235 2247
rect 1281 2201 1294 2247
rect 1222 2131 1294 2201
rect 1222 2085 1235 2131
rect 1281 2085 1294 2131
rect 1686 2317 1699 2363
rect 1745 2317 1758 2363
rect 1686 2247 1758 2317
rect 1686 2201 1699 2247
rect 1745 2201 1758 2247
rect 1686 2131 1758 2201
rect 1222 2028 1294 2085
rect 1686 2085 1699 2131
rect 1745 2085 1758 2131
rect 1686 2028 1758 2085
rect 1222 2015 1758 2028
rect 1222 1969 1235 2015
rect 1281 1969 1351 2015
rect 1397 1969 1467 2015
rect 1513 1969 1583 2015
rect 1629 1969 1699 2015
rect 1745 1969 1758 2015
rect 1222 1956 1758 1969
rect 73 1579 609 1592
rect 73 1533 86 1579
rect 132 1533 202 1579
rect 248 1533 318 1579
rect 364 1533 434 1579
rect 480 1533 550 1579
rect 596 1533 609 1579
rect 73 1520 609 1533
rect 73 1463 145 1520
rect 73 1417 86 1463
rect 132 1417 145 1463
rect 537 1463 609 1520
rect 73 1347 145 1417
rect 73 1301 86 1347
rect 132 1301 145 1347
rect 73 1231 145 1301
rect 73 1185 86 1231
rect 132 1185 145 1231
rect 537 1417 550 1463
rect 596 1417 609 1463
rect 537 1347 609 1417
rect 537 1301 550 1347
rect 596 1301 609 1347
rect 537 1231 609 1301
rect 73 1128 145 1185
rect 537 1185 550 1231
rect 596 1185 609 1231
rect 537 1128 609 1185
rect 73 1115 609 1128
rect 73 1069 86 1115
rect 132 1069 202 1115
rect 248 1069 318 1115
rect 364 1069 434 1115
rect 480 1069 550 1115
rect 596 1069 609 1115
rect 73 1056 609 1069
rect 1222 1579 1758 1592
rect 1222 1533 1235 1579
rect 1281 1533 1351 1579
rect 1397 1533 1467 1579
rect 1513 1533 1583 1579
rect 1629 1533 1699 1579
rect 1745 1533 1758 1579
rect 1222 1520 1758 1533
rect 1222 1463 1294 1520
rect 1222 1417 1235 1463
rect 1281 1417 1294 1463
rect 1686 1463 1758 1520
rect 1222 1347 1294 1417
rect 1222 1301 1235 1347
rect 1281 1301 1294 1347
rect 1222 1231 1294 1301
rect 1222 1185 1235 1231
rect 1281 1185 1294 1231
rect 1686 1417 1699 1463
rect 1745 1417 1758 1463
rect 1686 1347 1758 1417
rect 1686 1301 1699 1347
rect 1745 1301 1758 1347
rect 1686 1231 1758 1301
rect 1222 1128 1294 1185
rect 1686 1185 1699 1231
rect 1745 1185 1758 1231
rect 1686 1128 1758 1185
rect 1222 1115 1758 1128
rect 1222 1069 1235 1115
rect 1281 1069 1351 1115
rect 1397 1069 1467 1115
rect 1513 1069 1583 1115
rect 1629 1069 1699 1115
rect 1745 1069 1758 1115
rect 1222 1056 1758 1069
<< nsubdiffcont >>
rect 86 2433 132 2479
rect 202 2433 248 2479
rect 318 2433 364 2479
rect 434 2433 480 2479
rect 550 2433 596 2479
rect 86 2317 132 2363
rect 86 2201 132 2247
rect 86 2085 132 2131
rect 550 2317 596 2363
rect 550 2201 596 2247
rect 550 2085 596 2131
rect 86 1969 132 2015
rect 202 1969 248 2015
rect 318 1969 364 2015
rect 434 1969 480 2015
rect 550 1969 596 2015
rect 1235 2433 1281 2479
rect 1351 2433 1397 2479
rect 1467 2433 1513 2479
rect 1583 2433 1629 2479
rect 1699 2433 1745 2479
rect 1235 2317 1281 2363
rect 1235 2201 1281 2247
rect 1235 2085 1281 2131
rect 1699 2317 1745 2363
rect 1699 2201 1745 2247
rect 1699 2085 1745 2131
rect 1235 1969 1281 2015
rect 1351 1969 1397 2015
rect 1467 1969 1513 2015
rect 1583 1969 1629 2015
rect 1699 1969 1745 2015
rect 86 1533 132 1579
rect 202 1533 248 1579
rect 318 1533 364 1579
rect 434 1533 480 1579
rect 550 1533 596 1579
rect 86 1417 132 1463
rect 86 1301 132 1347
rect 86 1185 132 1231
rect 550 1417 596 1463
rect 550 1301 596 1347
rect 550 1185 596 1231
rect 86 1069 132 1115
rect 202 1069 248 1115
rect 318 1069 364 1115
rect 434 1069 480 1115
rect 550 1069 596 1115
rect 1235 1533 1281 1579
rect 1351 1533 1397 1579
rect 1467 1533 1513 1579
rect 1583 1533 1629 1579
rect 1699 1533 1745 1579
rect 1235 1417 1281 1463
rect 1235 1301 1281 1347
rect 1235 1185 1281 1231
rect 1699 1417 1745 1463
rect 1699 1301 1745 1347
rect 1699 1185 1745 1231
rect 1235 1069 1281 1115
rect 1351 1069 1397 1115
rect 1467 1069 1513 1115
rect 1583 1069 1629 1115
rect 1699 1069 1745 1115
<< pdiode >>
rect 241 2311 441 2324
rect 241 2265 254 2311
rect 300 2265 382 2311
rect 428 2265 441 2311
rect 241 2183 441 2265
rect 241 2137 254 2183
rect 300 2137 382 2183
rect 428 2137 441 2183
rect 241 2124 441 2137
rect 1390 2311 1590 2324
rect 1390 2265 1403 2311
rect 1449 2265 1531 2311
rect 1577 2265 1590 2311
rect 1390 2183 1590 2265
rect 1390 2137 1403 2183
rect 1449 2137 1531 2183
rect 1577 2137 1590 2183
rect 1390 2124 1590 2137
rect 241 1411 441 1424
rect 241 1365 254 1411
rect 300 1365 382 1411
rect 428 1365 441 1411
rect 241 1283 441 1365
rect 241 1237 254 1283
rect 300 1237 382 1283
rect 428 1237 441 1283
rect 241 1224 441 1237
rect 1390 1411 1590 1424
rect 1390 1365 1403 1411
rect 1449 1365 1531 1411
rect 1577 1365 1590 1411
rect 1390 1283 1590 1365
rect 1390 1237 1403 1283
rect 1449 1237 1531 1283
rect 1577 1237 1590 1283
rect 1390 1224 1590 1237
<< pdiodec >>
rect 254 2265 300 2311
rect 382 2265 428 2311
rect 254 2137 300 2183
rect 382 2137 428 2183
rect 1403 2265 1449 2311
rect 1531 2265 1577 2311
rect 1403 2137 1449 2183
rect 1531 2137 1577 2183
rect 254 1365 300 1411
rect 382 1365 428 1411
rect 254 1237 300 1283
rect 382 1237 428 1283
rect 1403 1365 1449 1411
rect 1531 1365 1577 1411
rect 1403 1237 1449 1283
rect 1531 1237 1577 1283
<< metal1 >>
rect 10095 7859 10347 7871
rect 10095 7703 10107 7859
rect 10159 7703 10347 7859
rect 10095 7691 10347 7703
rect 10275 7369 10351 7381
rect 10275 7213 10287 7369
rect 10339 7213 10351 7369
rect 10275 7201 10351 7213
rect 805 5974 881 5998
rect 805 5818 817 5974
rect 869 5873 881 5974
rect 1105 5987 1307 5998
rect 11632 5990 11688 6175
rect 1105 5935 1125 5987
rect 1281 5985 1307 5987
rect 11512 5985 11695 5990
rect 1281 5983 11695 5985
rect 1281 5935 11524 5983
rect 1105 5931 11524 5935
rect 11680 5931 11695 5983
rect 1105 5929 11695 5931
rect 1105 5924 1307 5929
rect 11512 5926 11695 5929
rect 12135 5901 12443 5902
rect 12738 5901 12986 6502
rect 11794 5873 11976 5877
rect 869 5871 11976 5873
rect 869 5819 11808 5871
rect 11964 5819 11976 5871
rect 869 5818 11976 5819
rect 805 5817 11976 5818
rect 805 5797 881 5817
rect 11794 5813 11976 5817
rect 12135 5853 12986 5901
rect 12135 5697 12158 5853
rect 12418 5697 12986 5853
rect 12135 5653 12986 5697
rect 12135 5652 12443 5653
rect 8310 5571 8815 5639
rect 9499 5571 9627 5639
rect 10570 5432 10873 5479
rect 10570 5380 10591 5432
rect 10851 5380 10873 5432
rect 10570 5335 10873 5380
rect 11170 5471 11265 5501
rect 11170 4691 11192 5471
rect 11244 5276 11265 5471
rect 13168 5362 13452 5374
rect 13168 5276 13388 5362
rect 11244 5109 13388 5276
rect 11244 4691 11265 5109
rect 13044 4894 13388 5109
rect 13440 4894 13452 5362
rect 13044 4882 13452 4894
rect 11170 4666 11265 4691
rect 377 4467 453 4479
rect 377 4311 389 4467
rect 441 4400 453 4467
rect 797 4467 873 4479
rect 797 4400 809 4467
rect 441 4311 809 4400
rect 861 4311 873 4467
rect 7991 4446 9118 4522
rect 13356 4458 13432 4470
rect 13356 4439 13368 4458
rect 12910 4326 13368 4439
rect 377 4299 873 4311
rect 13356 4302 13368 4326
rect 13420 4302 13432 4458
rect 13356 4290 13432 4302
rect 6820 4270 7000 4278
rect 6733 4266 7000 4270
rect 6733 4214 6832 4266
rect 6988 4214 7000 4266
rect 6733 4202 7000 4214
rect 11067 4076 11162 4104
rect 10629 3667 10841 3678
rect 2969 3347 3149 3359
rect 2969 3295 2981 3347
rect 3137 3295 3149 3347
rect 2969 3283 3149 3295
rect 10629 3303 10729 3667
rect 10781 3303 10841 3667
rect 10629 3292 10841 3303
rect 11067 3296 11083 4076
rect 11135 3755 11162 4076
rect 12136 3808 12316 3820
rect 12136 3756 12148 3808
rect 12304 3756 12316 3808
rect 12136 3755 12316 3756
rect 11135 3590 13041 3755
rect 11135 3296 11162 3590
rect 11067 3269 11162 3296
rect 7841 3169 9118 3245
rect 9499 3169 9627 3237
rect 3564 3078 5280 3090
rect 3564 3026 3581 3078
rect 3737 3026 5106 3078
rect 5262 3026 5280 3078
rect 3564 3013 5280 3026
rect 3171 2946 7115 2958
rect 3171 2894 3183 2946
rect 3339 2894 6943 2946
rect 7099 2894 7115 2946
rect 3171 2882 7115 2894
rect 9806 2669 11509 2681
rect -144 2625 2037 2637
rect -144 2573 -132 2625
rect 24 2573 2037 2625
rect 9806 2617 9818 2669
rect 9974 2617 11341 2669
rect 11497 2617 11509 2669
rect 9806 2605 11509 2617
rect -144 2561 2037 2573
rect 73 2479 609 2492
rect 73 2433 86 2479
rect 132 2433 202 2479
rect 248 2433 318 2479
rect 364 2433 434 2479
rect 480 2433 550 2479
rect 596 2433 609 2479
rect 73 2420 609 2433
rect 73 2363 145 2420
rect 73 2317 86 2363
rect 132 2317 145 2363
rect 537 2363 609 2420
rect 73 2247 145 2317
rect 73 2201 86 2247
rect 132 2201 145 2247
rect 73 2131 145 2201
rect 73 2085 86 2131
rect 132 2085 145 2131
rect 241 2311 441 2324
rect 241 2265 254 2311
rect 300 2265 382 2311
rect 428 2265 441 2311
rect 241 2250 441 2265
rect 241 2198 262 2250
rect 418 2198 441 2250
rect 241 2183 441 2198
rect 241 2137 254 2183
rect 300 2137 382 2183
rect 428 2137 441 2183
rect 241 2124 441 2137
rect 537 2317 550 2363
rect 596 2317 609 2363
rect 537 2247 609 2317
rect 537 2201 550 2247
rect 596 2201 609 2247
rect 537 2131 609 2201
rect 73 2028 145 2085
rect 537 2085 550 2131
rect 596 2085 609 2131
rect 537 2028 609 2085
rect 73 2015 609 2028
rect 73 1969 86 2015
rect 132 1969 202 2015
rect 248 1969 318 2015
rect 364 1969 434 2015
rect 480 1969 550 2015
rect 596 1969 609 2015
rect 73 1956 609 1969
rect 1222 2479 1758 2492
rect 1222 2433 1235 2479
rect 1281 2433 1351 2479
rect 1397 2433 1467 2479
rect 1513 2433 1583 2479
rect 1629 2433 1699 2479
rect 1745 2433 1758 2479
rect 1222 2420 1758 2433
rect 1222 2363 1294 2420
rect 1222 2317 1235 2363
rect 1281 2317 1294 2363
rect 1686 2363 1758 2420
rect 1222 2247 1294 2317
rect 1222 2201 1235 2247
rect 1281 2201 1294 2247
rect 1222 2131 1294 2201
rect 1222 2085 1235 2131
rect 1281 2085 1294 2131
rect 1390 2311 1590 2324
rect 1390 2265 1403 2311
rect 1449 2265 1531 2311
rect 1577 2265 1590 2311
rect 1390 2250 1590 2265
rect 1390 2198 1411 2250
rect 1567 2198 1590 2250
rect 1390 2183 1590 2198
rect 1390 2137 1403 2183
rect 1449 2137 1531 2183
rect 1577 2137 1590 2183
rect 1390 2124 1590 2137
rect 1686 2317 1699 2363
rect 1745 2317 1758 2363
rect 1686 2247 1758 2317
rect 1686 2201 1699 2247
rect 1745 2201 1758 2247
rect 1686 2131 1758 2201
rect 1222 2028 1294 2085
rect 1686 2085 1699 2131
rect 1745 2085 1758 2131
rect 1686 2028 1758 2085
rect 1961 2117 2037 2561
rect 2290 2361 3337 2566
rect 1961 2071 2351 2117
rect 2576 2071 2645 2117
rect 1222 2015 1758 2028
rect 1222 1969 1235 2015
rect 1281 1969 1351 2015
rect 1397 1969 1467 2015
rect 1513 1969 1583 2015
rect 1629 1969 1699 2015
rect 1745 1969 1758 2015
rect 1222 1956 1758 1969
rect 73 1713 1758 1956
rect 2533 1966 2585 1979
rect 2533 1797 2585 1810
rect 2826 1971 2879 1986
rect 2878 1815 2879 1971
rect 2826 1802 2879 1815
rect 73 1592 2975 1713
rect 73 1579 609 1592
rect 73 1533 86 1579
rect 132 1533 202 1579
rect 248 1533 318 1579
rect 364 1533 434 1579
rect 480 1533 550 1579
rect 596 1533 609 1579
rect 73 1520 609 1533
rect 73 1463 145 1520
rect 73 1417 86 1463
rect 132 1417 145 1463
rect 537 1463 609 1520
rect 73 1347 145 1417
rect 73 1301 86 1347
rect 132 1301 145 1347
rect 73 1231 145 1301
rect 73 1185 86 1231
rect 132 1185 145 1231
rect 241 1411 441 1424
rect 241 1403 254 1411
rect 300 1403 382 1411
rect 241 1247 253 1403
rect 305 1365 382 1403
rect 428 1365 441 1411
rect 305 1283 441 1365
rect 305 1247 382 1283
rect 241 1237 254 1247
rect 300 1237 382 1247
rect 428 1237 441 1283
rect 241 1224 441 1237
rect 537 1417 550 1463
rect 596 1417 609 1463
rect 537 1347 609 1417
rect 537 1301 550 1347
rect 596 1301 609 1347
rect 537 1231 609 1301
rect 73 1128 145 1185
rect 537 1185 550 1231
rect 596 1185 609 1231
rect 537 1128 609 1185
rect 73 1115 609 1128
rect 73 1069 86 1115
rect 132 1069 202 1115
rect 248 1069 318 1115
rect 364 1069 434 1115
rect 480 1069 550 1115
rect 596 1069 609 1115
rect 73 1056 609 1069
rect 1222 1579 2975 1592
rect 1222 1533 1235 1579
rect 1281 1533 1351 1579
rect 1397 1533 1467 1579
rect 1513 1533 1583 1579
rect 1629 1533 1699 1579
rect 1745 1540 2975 1579
rect 1745 1533 1758 1540
rect 1222 1520 1758 1533
rect 1222 1463 1294 1520
rect 1222 1417 1235 1463
rect 1281 1417 1294 1463
rect 1686 1463 1758 1520
rect 1222 1347 1294 1417
rect 1222 1301 1235 1347
rect 1281 1301 1294 1347
rect 1222 1231 1294 1301
rect 1222 1185 1235 1231
rect 1281 1185 1294 1231
rect 1390 1411 1590 1424
rect 1390 1365 1403 1411
rect 1449 1365 1531 1411
rect 1577 1365 1590 1411
rect 1390 1350 1590 1365
rect 1390 1298 1411 1350
rect 1567 1298 1590 1350
rect 1390 1283 1590 1298
rect 1390 1237 1403 1283
rect 1449 1237 1531 1283
rect 1577 1237 1590 1283
rect 1390 1224 1590 1237
rect 1686 1417 1699 1463
rect 1745 1417 1758 1463
rect 1686 1347 1758 1417
rect 1686 1301 1699 1347
rect 1745 1301 1758 1347
rect 1686 1231 1758 1301
rect 1222 1128 1294 1185
rect 1686 1185 1699 1231
rect 1745 1185 1758 1231
rect 1686 1128 1758 1185
rect 1222 1115 1758 1128
rect 1222 1069 1235 1115
rect 1281 1069 1351 1115
rect 1397 1069 1467 1115
rect 1513 1069 1583 1115
rect 1629 1069 1699 1115
rect 1745 1069 1758 1115
rect 1222 1056 1758 1069
rect 73 939 2971 1056
rect 73 893 2306 939
rect 2352 893 2599 939
rect 2645 893 2892 939
rect 2938 893 2971 939
rect 73 886 2971 893
rect 73 686 1843 886
rect 2535 769 2587 781
rect 73 683 1833 686
rect 2043 611 2119 623
rect 2043 455 2055 611
rect 2107 516 2119 611
rect 2535 601 2587 613
rect 2829 774 2881 786
rect 2829 606 2881 618
rect 2107 470 2351 516
rect 2580 470 2642 516
rect 2107 455 2119 470
rect 2043 444 2119 455
rect 3132 235 3337 2361
rect 11406 2125 11482 2138
rect 11406 1969 11418 2125
rect 11470 1969 11482 2125
rect 11406 1956 11482 1969
rect 7988 1465 8218 1474
rect 7988 1413 8025 1465
rect 8181 1413 8218 1465
rect 7988 1405 8218 1413
rect 8463 1464 8693 1473
rect 8463 1412 8500 1464
rect 8656 1412 8693 1464
rect 8463 1404 8693 1412
rect 12366 1464 12596 1473
rect 12366 1412 12403 1464
rect 12559 1412 12596 1464
rect 12366 1404 12596 1412
rect 4077 1377 4339 1400
rect 4077 1325 4126 1377
rect 4282 1325 4339 1377
rect 4077 1303 4339 1325
rect 4091 1173 4321 1182
rect 4091 1121 4128 1173
rect 4284 1121 4321 1173
rect 7986 1181 8216 1190
rect 7986 1129 8023 1181
rect 8179 1129 8216 1181
rect 7986 1121 8216 1129
rect 8465 1180 8695 1189
rect 8465 1128 8502 1180
rect 8658 1128 8695 1180
rect 4091 1113 4321 1121
rect 8465 1120 8695 1128
rect 12364 1180 12594 1189
rect 12364 1128 12401 1180
rect 12557 1128 12594 1180
rect 12364 1120 12594 1128
rect 2293 30 3337 235
<< via1 >>
rect 10107 7703 10159 7859
rect 10287 7213 10339 7369
rect 817 5818 869 5974
rect 1125 5935 1281 5987
rect 11524 5931 11680 5983
rect 11808 5819 11964 5871
rect 12158 5697 12418 5853
rect 10591 5380 10851 5432
rect 11192 4691 11244 5471
rect 13388 4894 13440 5362
rect 389 4311 441 4467
rect 809 4311 861 4467
rect 13368 4302 13420 4458
rect 6832 4214 6988 4266
rect 2981 3295 3137 3347
rect 10729 3303 10781 3667
rect 11083 3296 11135 4076
rect 12148 3756 12304 3808
rect 3581 3026 3737 3078
rect 5106 3026 5262 3078
rect 3183 2894 3339 2946
rect 6943 2894 7099 2946
rect -132 2573 24 2625
rect 9818 2617 9974 2669
rect 11341 2617 11497 2669
rect 262 2198 418 2250
rect 1411 2198 1567 2250
rect 2533 1810 2585 1966
rect 2826 1815 2878 1971
rect 253 1365 254 1403
rect 254 1365 300 1403
rect 300 1365 305 1403
rect 253 1283 305 1365
rect 253 1247 254 1283
rect 254 1247 300 1283
rect 300 1247 305 1283
rect 1411 1298 1567 1350
rect 2055 455 2107 611
rect 2535 613 2587 769
rect 2829 618 2881 774
rect 5216 1967 5268 2123
rect 7044 1968 7096 2124
rect 10078 1969 10130 2125
rect 11418 1969 11470 2125
rect 8025 1413 8181 1465
rect 8500 1412 8656 1464
rect 12403 1412 12559 1464
rect 4126 1325 4282 1377
rect 4128 1121 4284 1173
rect 8023 1129 8179 1181
rect 8502 1128 8658 1180
rect 12401 1128 12557 1180
<< metal2 >>
rect 10095 7859 10171 7871
rect 10095 7703 10107 7859
rect 10159 7703 10171 7859
rect 10095 6313 10171 7703
rect 805 5974 881 5998
rect 805 5818 817 5974
rect 869 5818 881 5974
rect 1106 5987 1307 5998
rect 1106 5935 1125 5987
rect 1281 5935 1307 5987
rect 1106 5924 1307 5935
rect 805 5797 881 5818
rect 805 4479 869 5797
rect 377 4467 453 4479
rect 377 4311 389 4467
rect 441 4311 453 4467
rect -144 2625 36 2637
rect -144 2573 -132 2625
rect 24 2573 36 2625
rect -144 2561 36 2573
rect -144 1415 -68 2561
rect 377 2262 453 4311
rect 797 4467 873 4479
rect 797 4311 809 4467
rect 861 4311 873 4467
rect 1108 4393 1172 5924
rect 6579 5511 6779 6291
rect 9910 6237 10171 6313
rect 10275 7369 10351 7381
rect 10275 7213 10287 7369
rect 10339 7213 10351 7369
rect 6579 5351 7000 5511
rect 1108 4317 1328 4393
rect 797 4299 873 4311
rect 250 2250 453 2262
rect 250 2198 262 2250
rect 418 2198 453 2250
rect 250 2186 453 2198
rect 1252 2262 1328 4317
rect 6820 4266 7000 4278
rect 6820 4214 6832 4266
rect 6988 4214 7000 4266
rect 6820 4202 7000 4214
rect 2295 3129 2371 4152
rect 2969 3348 3149 3359
rect 2969 3347 3640 3348
rect 2969 3295 2981 3347
rect 3137 3295 3640 3347
rect 2969 3272 3640 3295
rect 2295 3053 3237 3129
rect 3161 2958 3237 3053
rect 3564 3090 3640 3272
rect 3564 3078 3752 3090
rect 3564 3026 3581 3078
rect 3737 3026 3752 3078
rect 3564 3013 3752 3026
rect 5093 3078 5280 3090
rect 5093 3026 5106 3078
rect 5262 3026 5280 3078
rect 5093 3013 5280 3026
rect 3161 2946 3351 2958
rect 3161 2894 3183 2946
rect 3339 2894 3351 2946
rect 3161 2882 3351 2894
rect 1252 2250 1589 2262
rect 1252 2198 1411 2250
rect 1567 2198 1589 2250
rect 1252 2186 1589 2198
rect -144 1403 317 1415
rect -144 1247 253 1403
rect 305 1247 317 1403
rect -144 1235 317 1247
rect -144 422 -68 1235
rect 377 422 453 2186
rect 2520 2071 3071 2133
rect 2520 1980 2582 2071
rect 2520 1966 2590 1980
rect 2520 1810 2533 1966
rect 2585 1810 2590 1966
rect 2520 1778 2590 1810
rect 2820 1971 2882 1985
rect 2820 1815 2826 1971
rect 2878 1815 2882 1971
rect 2520 1771 2582 1778
rect 2820 1603 2882 1815
rect 3009 1665 3071 2071
rect 5204 2123 5280 3013
rect 6931 2946 7115 2958
rect 6931 2894 6943 2946
rect 7099 2894 7115 2946
rect 6931 2882 7115 2894
rect 5204 1967 5216 2123
rect 5268 1967 5280 2123
rect 5204 1954 5280 1967
rect 7033 2124 7108 2882
rect 9910 2681 9986 6237
rect 10275 6177 10351 7213
rect 9806 2669 9986 2681
rect 9806 2617 9818 2669
rect 9974 2617 9986 2669
rect 9806 2605 9986 2617
rect 10066 6100 10351 6177
rect 7033 1968 7044 2124
rect 7096 1968 7108 2124
rect 7033 1952 7108 1968
rect 10066 2125 10142 6100
rect 11130 5637 11186 6529
rect 11282 5765 11338 6529
rect 11632 5990 11688 6175
rect 11512 5983 11695 5990
rect 11512 5931 11524 5983
rect 11680 5931 11695 5983
rect 11512 5926 11695 5931
rect 11907 5877 11963 6369
rect 11794 5871 11976 5877
rect 11794 5819 11808 5871
rect 11964 5819 11976 5871
rect 11794 5813 11976 5819
rect 12135 5853 12443 5902
rect 11282 5709 11538 5765
rect 11130 5581 11386 5637
rect 11170 5479 11265 5501
rect 10570 5471 11265 5479
rect 10570 5432 11192 5471
rect 10570 5380 10591 5432
rect 10851 5380 11192 5432
rect 10570 5335 11192 5380
rect 11170 4691 11192 5335
rect 11244 4691 11265 5471
rect 11170 4666 11265 4691
rect 11067 4076 11162 4104
rect 11067 3678 11083 4076
rect 10670 3667 11083 3678
rect 10670 3303 10729 3667
rect 10781 3303 11083 3667
rect 10670 3296 11083 3303
rect 11135 3296 11162 4076
rect 10670 3292 11162 3296
rect 11067 3269 11162 3292
rect 11330 3049 11386 5581
rect 10066 1969 10078 2125
rect 10130 1969 10142 2125
rect 10066 1954 10142 1969
rect 10858 2992 11386 3049
rect 3009 1645 5902 1665
rect 3009 1603 8016 1645
rect 2817 1546 2882 1603
rect 5840 1583 8016 1603
rect 2820 1528 2882 1546
rect 2820 1508 5768 1528
rect 2820 1466 7833 1508
rect 7954 1488 8016 1583
rect 5706 1446 7833 1466
rect 4077 1377 4358 1400
rect 4077 1375 4126 1377
rect 1399 1350 2119 1362
rect 1399 1298 1411 1350
rect 1567 1298 2119 1350
rect 1399 1286 2119 1298
rect 2043 611 2119 1286
rect 3904 1325 4126 1375
rect 4282 1325 4358 1377
rect 3904 1313 4358 1325
rect 3904 1254 3966 1313
rect 4077 1303 4358 1313
rect 2043 455 2055 611
rect 2107 455 2119 611
rect 2530 1192 3966 1254
rect 2530 769 2592 1192
rect 4075 1173 4356 1200
rect 4075 1122 4128 1173
rect 2530 613 2535 769
rect 2587 613 2592 769
rect 2530 599 2592 613
rect 2823 1121 4128 1122
rect 4284 1121 4356 1173
rect 7772 1198 7833 1446
rect 7949 1465 8230 1488
rect 7949 1413 8025 1465
rect 8181 1413 8230 1465
rect 7949 1391 8230 1413
rect 8451 1464 8732 1487
rect 8451 1412 8500 1464
rect 8656 1412 9005 1464
rect 8451 1407 9005 1412
rect 8451 1390 8732 1407
rect 8948 1367 9005 1407
rect 10858 1367 10915 2992
rect 11482 2930 11538 5709
rect 12135 5697 12158 5853
rect 12418 5697 12443 5853
rect 12135 5652 12443 5697
rect 12136 3808 12316 5652
rect 12136 3756 12148 3808
rect 12304 3756 12316 3808
rect 12136 3348 12316 3756
rect 12136 3292 12146 3348
rect 12306 3292 12316 3348
rect 12136 3278 12316 3292
rect 8948 1310 10915 1367
rect 10982 2874 11538 2930
rect 10982 1240 11038 2874
rect 11329 2669 11509 2681
rect 11329 2617 11341 2669
rect 11497 2617 11509 2669
rect 11329 2605 11509 2617
rect 11406 2125 11482 2605
rect 11406 1969 11418 2125
rect 11470 1969 11482 2125
rect 11406 1956 11482 1969
rect 12528 1487 12584 6511
rect 12660 2820 12716 6511
rect 13376 5364 13452 5374
rect 13376 4892 13386 5364
rect 13442 4892 13452 5364
rect 13376 4882 13452 4892
rect 13356 4458 13432 4470
rect 13356 4302 13368 4458
rect 13420 4302 13432 4458
rect 13356 4290 13432 4302
rect 12660 2741 12726 2820
rect 12327 1464 12608 1487
rect 12327 1412 12403 1464
rect 12559 1412 12608 1464
rect 12327 1390 12608 1412
rect 7951 1198 8232 1208
rect 7772 1181 8232 1198
rect 7772 1137 8023 1181
rect 2823 1103 4356 1121
rect 7951 1129 8023 1137
rect 8179 1129 8232 1181
rect 7951 1111 8232 1129
rect 8449 1181 8730 1207
rect 8972 1184 11038 1240
rect 8972 1181 9028 1184
rect 8449 1180 9028 1181
rect 8449 1128 8502 1180
rect 8658 1128 9028 1180
rect 8449 1125 9028 1128
rect 12329 1180 12610 1207
rect 12329 1128 12401 1180
rect 12557 1169 12610 1180
rect 12670 1169 12726 2741
rect 12557 1128 12726 1169
rect 8449 1110 8730 1125
rect 12329 1113 12726 1128
rect 12329 1110 12610 1113
rect 2823 1060 4171 1103
rect 2823 774 2885 1060
rect 2823 618 2829 774
rect 2881 618 2885 774
rect 2823 601 2885 618
rect 2043 444 2119 455
<< via2 >>
rect 12146 3292 12306 3348
rect 13386 5362 13442 5364
rect 13386 4894 13388 5362
rect 13388 4894 13440 5362
rect 13440 4894 13442 5362
rect 13386 4892 13442 4894
<< metal3 >>
rect 9619 4882 9695 5374
rect 13376 5364 13452 5374
rect 13376 4892 13386 5364
rect 13442 4892 13452 5364
rect 13376 4882 13452 4892
rect 9619 3696 9695 4188
rect 12136 3348 12316 3358
rect 12136 3292 12146 3348
rect 12306 3292 12316 3348
rect 12136 3282 12316 3292
use comp018green_in_cms_smt  comp018green_in_cms_smt_0
timestamp 1764353313
transform 1 0 1532 0 1 3158
box -1470 -83 6875 2578
use comp018green_in_drv  comp018green_in_drv_0
timestamp 1764353313
transform 1 0 8900 0 1 3158
box -496 -83 4246 2578
use comp018green_in_logic_pupd  comp018green_in_logic_pupd_0
timestamp 1764353313
transform -1 0 13932 0 1 9724
box 946 -3664 2905 1086
use comp018green_in_pupd  comp018green_in_pupd_0
timestamp 1764353313
transform 0 -1 2979 -1 0 14857
box -83 -7815 8792 3035
use comp018green_sigbuf  comp018green_sigbuf_0
timestamp 1764353313
transform 1 0 7863 0 -1 2492
box 349 -83 2798 2578
use comp018green_sigbuf  comp018green_sigbuf_1
timestamp 1764353313
transform 1 0 3489 0 -1 2492
box 349 -83 2798 2578
use comp018green_sigbuf  comp018green_sigbuf_2
timestamp 1764353313
transform -1 0 13197 0 -1 2492
box 349 -83 2798 2578
use comp018green_sigbuf  comp018green_sigbuf_3
timestamp 1764353313
transform -1 0 8823 0 -1 2492
box 349 -83 2798 2578
use lv_inv  lv_inv_14
timestamp 1764353313
transform 1 0 -13774 0 1 -50649
box 15980 50799 16518 51697
use lv_inv  lv_inv_15
timestamp 1764353313
transform 1 0 -13480 0 1 -50649
box 15980 50799 16518 51697
use lv_inv  lv_inv_18
timestamp 1764353313
transform 1 0 -13776 0 -1 53236
box 15980 50799 16518 51697
use lv_inv  lv_inv_19
timestamp 1764353313
transform 1 0 -13482 0 -1 53236
box 15980 50799 16518 51697
<< labels >>
rlabel metal2 s 6679 6191 6679 6191 4 PAD
port 1 nsew
rlabel metal2 s -107 526 -107 526 4 CS
port 2 nsew
rlabel metal2 s 414 522 414 522 4 PU
port 3 nsew
<< properties >>
string GDS_END 10708276
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 10677192
<< end >>
