magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect 16870 51136 17574 51686
<< nmos >>
rect 17148 50930 17204 51050
rect 17280 50930 17336 51050
<< pmos >>
rect 17113 51222 17169 51462
rect 17280 51222 17336 51462
<< ndiff >>
rect 17059 51014 17148 51050
rect 17059 50968 17073 51014
rect 17119 50968 17148 51014
rect 17059 50930 17148 50968
rect 17204 50930 17280 51050
rect 17336 51013 17424 51050
rect 17336 50967 17365 51013
rect 17411 50967 17424 51013
rect 17336 50930 17424 50967
<< pdiff >>
rect 17024 51412 17113 51462
rect 17024 51272 17038 51412
rect 17084 51272 17113 51412
rect 17024 51222 17113 51272
rect 17169 51404 17280 51462
rect 17169 51358 17200 51404
rect 17246 51358 17280 51404
rect 17169 51222 17280 51358
rect 17336 51411 17424 51462
rect 17336 51271 17365 51411
rect 17411 51271 17424 51411
rect 17336 51222 17424 51271
<< ndiffc >>
rect 17073 50968 17119 51014
rect 17365 50967 17411 51013
<< pdiffc >>
rect 17038 51272 17084 51412
rect 17200 51358 17246 51404
rect 17365 51271 17411 51411
<< psubdiff >>
rect 16960 50849 17488 50864
rect 16960 50803 16973 50849
rect 17019 50803 17429 50849
rect 17475 50803 17488 50849
rect 16960 50788 17488 50803
<< nsubdiff >>
rect 16956 51589 17488 51604
rect 16956 51543 16973 51589
rect 17019 51543 17429 51589
rect 17475 51543 17488 51589
rect 16956 51528 17488 51543
<< psubdiffcont >>
rect 16973 50803 17019 50849
rect 17429 50803 17475 50849
<< nsubdiffcont >>
rect 16973 51543 17019 51589
rect 17429 51543 17475 51589
<< polysilicon >>
rect 17113 51462 17169 51506
rect 17280 51462 17336 51506
rect 17113 51168 17169 51222
rect 17113 51154 17204 51168
rect 17280 51167 17336 51222
rect 17113 51108 17134 51154
rect 17180 51108 17204 51154
rect 17113 51095 17204 51108
rect 17252 51154 17336 51167
rect 17252 51108 17270 51154
rect 17316 51108 17336 51154
rect 17252 51095 17336 51108
rect 17148 51050 17204 51095
rect 17280 51050 17336 51095
rect 17148 50885 17204 50930
rect 17280 50886 17336 50930
<< polycontact >>
rect 17134 51108 17180 51154
rect 17270 51108 17316 51154
<< metal1 >>
rect 16956 51589 17488 51600
rect 16956 51543 16973 51589
rect 17019 51543 17429 51589
rect 17475 51543 17488 51589
rect 16956 51525 17488 51543
rect 17038 51412 17084 51461
rect 17179 51404 17270 51525
rect 17179 51358 17200 51404
rect 17246 51358 17270 51404
rect 17179 51304 17270 51358
rect 17365 51411 17411 51459
rect 17038 51258 17084 51272
rect 17365 51258 17411 51271
rect 17038 51211 17411 51258
rect 17059 51154 17218 51165
rect 17059 51108 17134 51154
rect 17180 51108 17218 51154
rect 17059 51094 17218 51108
rect 17268 51154 17318 51165
rect 17268 51108 17270 51154
rect 17316 51108 17318 51154
rect 17073 51014 17119 51048
rect 17268 51046 17318 51108
rect 17073 50868 17119 50968
rect 17213 50983 17318 51046
rect 17365 51013 17411 51211
rect 17213 50940 17271 50983
rect 17365 50933 17411 50967
rect 16960 50849 17488 50868
rect 16960 50803 16973 50849
rect 17019 50803 17429 50849
rect 17475 50803 17488 50849
rect 16960 50792 17488 50803
<< properties >>
string GDS_END 10537418
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 10534534
<< end >>
