magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect -5 111 12385 13626
<< psubdiff >>
rect -767 15239 13147 15294
rect -767 14593 -745 15239
rect 901 14593 1299 15239
rect -767 14481 1299 14593
rect -767 -865 -733 14481
rect -87 13693 1299 14481
rect 2245 13693 3071 15239
rect 4017 13693 4836 15239
rect 5782 13693 6605 15239
rect 7551 13693 8374 15239
rect 9320 13693 10140 15239
rect 11086 15234 13147 15239
rect 11086 14588 11479 15234
rect 13125 14588 13147 15234
rect 11086 14481 13147 14588
rect 11086 13693 12467 14481
rect -87 13666 12467 13693
rect -87 63 -53 13666
rect 12433 63 12467 13666
rect -87 41 12467 63
rect -87 -805 118 41
rect 12264 -805 12467 41
rect -87 -865 12467 -805
rect 13113 -865 13147 14481
rect -767 -938 13147 -865
rect -767 -1284 -733 -938
rect 13113 -1284 13147 -938
rect -767 -1312 13147 -1284
<< nsubdiff >>
rect 81 13500 12299 13540
rect 81 13479 1318 13500
rect 81 13133 103 13479
rect 849 13133 1318 13479
rect 81 12990 1318 13133
rect 81 1100 159 12990
rect 393 12958 1318 12990
rect 393 11596 624 12958
rect 858 11596 1318 12958
rect 393 11554 1318 11596
rect 2264 11554 3018 13500
rect 4064 11554 4818 13500
rect 5764 11554 6618 13500
rect 7564 11554 8318 13500
rect 9364 11554 10118 13500
rect 11064 13479 12299 13500
rect 11064 13133 11531 13479
rect 12277 13133 12299 13479
rect 11064 12990 12299 13133
rect 11064 12958 11987 12990
rect 11064 11596 11524 12958
rect 11758 11596 11987 12958
rect 11064 11554 11987 11596
rect 393 11504 11987 11554
rect 393 2431 451 11504
rect 11931 2431 11987 11504
rect 393 2409 11987 2431
rect 393 1163 636 2409
rect 11782 1163 11987 2409
rect 393 1100 11987 1163
rect 12221 1100 12299 12990
rect 81 1014 12299 1100
rect 81 268 118 1014
rect 12264 268 12299 1014
rect 81 246 12299 268
<< psubdiffcont >>
rect -745 14593 901 15239
rect -733 -865 -87 14481
rect 1299 13693 2245 15239
rect 3071 13693 4017 15239
rect 4836 13693 5782 15239
rect 6605 13693 7551 15239
rect 8374 13693 9320 15239
rect 10140 13693 11086 15239
rect 11479 14588 13125 15234
rect 118 -805 12264 41
rect 12467 -865 13113 14481
rect -733 -1284 13113 -938
<< nsubdiffcont >>
rect 103 13133 849 13479
rect 159 1100 393 12990
rect 624 11596 858 12958
rect 1318 11554 2264 13500
rect 3018 11554 4064 13500
rect 4818 11554 5764 13500
rect 6618 11554 7564 13500
rect 8318 11554 9364 13500
rect 10118 11554 11064 13500
rect 11531 13133 12277 13479
rect 11524 11596 11758 12958
rect 636 1163 11782 2409
rect 11987 1100 12221 12990
rect 118 268 12264 1014
<< polysilicon >>
rect 974 11125 1185 11144
rect 974 11079 1009 11125
rect 1149 11079 1185 11125
rect 974 11060 1185 11079
rect 2360 11125 2571 11144
rect 2360 11079 2395 11125
rect 2535 11079 2571 11125
rect 2360 11060 2571 11079
rect 2746 11125 2957 11144
rect 2746 11079 2781 11125
rect 2921 11079 2957 11125
rect 2746 11060 2957 11079
rect 4120 11125 4331 11144
rect 4120 11079 4155 11125
rect 4295 11079 4331 11125
rect 4120 11060 4331 11079
rect 4511 11125 4722 11144
rect 4511 11079 4546 11125
rect 4686 11079 4722 11125
rect 4511 11060 4722 11079
rect 5892 11125 6103 11144
rect 5892 11079 5927 11125
rect 6067 11079 6103 11125
rect 5892 11060 6103 11079
rect 6280 11125 6491 11144
rect 6280 11079 6315 11125
rect 6455 11079 6491 11125
rect 6280 11060 6491 11079
rect 7662 11125 7873 11144
rect 7662 11079 7697 11125
rect 7837 11079 7873 11125
rect 7662 11060 7873 11079
rect 8049 11125 8260 11144
rect 8049 11079 8084 11125
rect 8224 11079 8260 11125
rect 8049 11060 8260 11079
rect 9428 11125 9639 11144
rect 9428 11079 9463 11125
rect 9603 11079 9639 11125
rect 9428 11060 9639 11079
rect 9815 11125 10026 11144
rect 9815 11079 9850 11125
rect 9990 11079 10026 11125
rect 9815 11060 10026 11079
rect 11201 11125 11412 11144
rect 11201 11079 11236 11125
rect 11376 11079 11412 11125
rect 11201 11060 11412 11079
rect 974 2865 1185 2884
rect 974 2819 1009 2865
rect 1149 2819 1185 2865
rect 974 2800 1185 2819
rect 2360 2865 2571 2884
rect 2360 2819 2395 2865
rect 2535 2819 2571 2865
rect 2360 2800 2571 2819
rect 2746 2865 2957 2884
rect 2746 2819 2781 2865
rect 2921 2819 2957 2865
rect 2746 2800 2957 2819
rect 4120 2865 4331 2884
rect 4120 2819 4155 2865
rect 4295 2819 4331 2865
rect 4120 2800 4331 2819
rect 4511 2865 4722 2884
rect 4511 2819 4546 2865
rect 4686 2819 4722 2865
rect 4511 2800 4722 2819
rect 5892 2865 6103 2884
rect 5892 2819 5927 2865
rect 6067 2819 6103 2865
rect 5892 2800 6103 2819
rect 6280 2865 6491 2884
rect 6280 2819 6315 2865
rect 6455 2819 6491 2865
rect 6280 2800 6491 2819
rect 7662 2865 7873 2884
rect 7662 2819 7697 2865
rect 7837 2819 7873 2865
rect 7662 2800 7873 2819
rect 8049 2865 8260 2884
rect 8049 2819 8084 2865
rect 8224 2819 8260 2865
rect 8049 2800 8260 2819
rect 9428 2865 9639 2884
rect 9428 2819 9463 2865
rect 9603 2819 9639 2865
rect 9428 2800 9639 2819
rect 9815 2865 10026 2884
rect 9815 2819 9850 2865
rect 9990 2819 10026 2865
rect 9815 2800 10026 2819
rect 11201 2865 11412 2884
rect 11201 2819 11236 2865
rect 11376 2819 11412 2865
rect 11201 2800 11412 2819
<< polycontact >>
rect 1009 11079 1149 11125
rect 2395 11079 2535 11125
rect 2781 11079 2921 11125
rect 4155 11079 4295 11125
rect 4546 11079 4686 11125
rect 5927 11079 6067 11125
rect 6315 11079 6455 11125
rect 7697 11079 7837 11125
rect 8084 11079 8224 11125
rect 9463 11079 9603 11125
rect 9850 11079 9990 11125
rect 11236 11079 11376 11125
rect 1009 2819 1149 2865
rect 2395 2819 2535 2865
rect 2781 2819 2921 2865
rect 4155 2819 4295 2865
rect 4546 2819 4686 2865
rect 5927 2819 6067 2865
rect 6315 2819 6455 2865
rect 7697 2819 7837 2865
rect 8084 2819 8224 2865
rect 9463 2819 9603 2865
rect 9850 2819 9990 2865
rect 11236 2819 11376 2865
<< metal1 >>
rect -756 15239 912 15250
rect -756 14593 -745 15239
rect 901 14593 912 15239
rect -756 14548 -719 14593
rect -667 14548 -611 14593
rect -559 14548 -503 14593
rect -451 14582 912 14593
rect 1288 15239 2256 15250
rect -451 14548 -64 14582
rect -756 14492 -64 14548
rect -756 14481 -719 14492
rect -667 14481 -611 14492
rect -559 14481 -503 14492
rect -451 14481 -64 14492
rect -756 -865 -733 14481
rect -87 52 -64 14481
rect 1288 13693 1299 15239
rect 2245 13693 2256 15239
rect 1288 13682 2256 13693
rect 3060 15239 4028 15250
rect 3060 13693 3071 15239
rect 4017 13693 4028 15239
rect 3060 13682 4028 13693
rect 4825 15239 5793 15250
rect 4825 13693 4836 15239
rect 5782 13693 5793 15239
rect 4825 13682 5793 13693
rect 6594 15239 7562 15250
rect 6594 13693 6605 15239
rect 7551 13693 7562 15239
rect 6594 13682 7562 13693
rect 8363 15239 9331 15250
rect 8363 13693 8374 15239
rect 9320 13693 9331 15239
rect 8363 13682 9331 13693
rect 10129 15239 11097 15250
rect 10129 13693 10140 15239
rect 11086 13693 11097 15239
rect 11468 15234 13136 15245
rect 11468 14588 11479 15234
rect 13125 14588 13136 15234
rect 11468 14577 13136 14588
rect 10129 13682 11097 13693
rect 12444 14481 13136 14577
rect 1267 13500 2286 13540
rect 92 13479 889 13490
rect 92 13133 103 13479
rect 849 13133 889 13479
rect 92 13109 889 13133
rect 92 13057 472 13109
rect 524 13057 596 13109
rect 648 13057 720 13109
rect 772 13057 889 13109
rect 92 13029 889 13057
rect 142 12990 889 13029
rect 142 1100 159 12990
rect 393 12985 889 12990
rect 393 12933 472 12985
rect 524 12933 596 12985
rect 648 12958 720 12985
rect 772 12958 889 12985
rect 393 12861 624 12933
rect 393 12809 472 12861
rect 524 12809 596 12861
rect 393 12737 624 12809
rect 393 12685 472 12737
rect 524 12685 596 12737
rect 393 12613 624 12685
rect 393 12561 472 12613
rect 524 12561 596 12613
rect 393 12489 624 12561
rect 393 12437 472 12489
rect 524 12437 596 12489
rect 393 12365 624 12437
rect 393 12313 472 12365
rect 524 12313 596 12365
rect 393 12241 624 12313
rect 393 12189 472 12241
rect 524 12189 596 12241
rect 393 12117 624 12189
rect 393 12065 472 12117
rect 524 12065 596 12117
rect 393 11993 624 12065
rect 393 11941 472 11993
rect 524 11941 596 11993
rect 393 11869 624 11941
rect 393 11817 472 11869
rect 524 11817 596 11869
rect 393 11745 624 11817
rect 393 11693 472 11745
rect 524 11693 596 11745
rect 393 11621 624 11693
rect 393 11569 472 11621
rect 524 11569 596 11621
rect 858 11596 889 12958
rect 648 11569 720 11596
rect 772 11569 889 11596
rect 393 11543 889 11569
rect 1267 11554 1318 13500
rect 2264 11554 2286 13500
rect 1267 11543 2286 11554
rect 2983 13500 4093 13540
rect 2983 11554 3018 13500
rect 4064 11554 4093 13500
rect 2983 11543 4093 11554
rect 4768 13500 5799 13540
rect 4768 11554 4818 13500
rect 5764 11554 5799 13500
rect 4768 11543 5799 11554
rect 6570 13500 7605 13540
rect 6570 11554 6618 13500
rect 7564 11554 7605 13500
rect 6570 11543 7605 11554
rect 8286 13500 9398 13540
rect 8286 11554 8318 13500
rect 9364 11554 9398 13500
rect 8286 11543 9398 11554
rect 10079 13500 11105 13540
rect 10079 11554 10118 13500
rect 11064 11554 11105 13500
rect 10079 11543 11105 11554
rect 11498 13479 12288 13490
rect 11498 13133 11531 13479
rect 12277 13133 12288 13479
rect 11498 13109 12288 13133
rect 11498 13057 11601 13109
rect 11653 13057 11725 13109
rect 11777 13057 11849 13109
rect 11901 13057 12288 13109
rect 11498 13029 12288 13057
rect 11498 12990 12238 13029
rect 11498 12985 11987 12990
rect 11498 12958 11601 12985
rect 11653 12958 11725 12985
rect 11498 11596 11524 12958
rect 11777 12933 11849 12985
rect 11901 12933 11987 12985
rect 11758 12861 11987 12933
rect 11777 12809 11849 12861
rect 11901 12809 11987 12861
rect 11758 12737 11987 12809
rect 11777 12685 11849 12737
rect 11901 12685 11987 12737
rect 11758 12613 11987 12685
rect 11777 12561 11849 12613
rect 11901 12561 11987 12613
rect 11758 12489 11987 12561
rect 11777 12437 11849 12489
rect 11901 12437 11987 12489
rect 11758 12365 11987 12437
rect 11777 12313 11849 12365
rect 11901 12313 11987 12365
rect 11758 12241 11987 12313
rect 11777 12189 11849 12241
rect 11901 12189 11987 12241
rect 11758 12117 11987 12189
rect 11777 12065 11849 12117
rect 11901 12065 11987 12117
rect 11758 11993 11987 12065
rect 11777 11941 11849 11993
rect 11901 11941 11987 11993
rect 11758 11869 11987 11941
rect 11777 11817 11849 11869
rect 11901 11817 11987 11869
rect 11758 11745 11987 11817
rect 11777 11693 11849 11745
rect 11901 11693 11987 11745
rect 11758 11621 11987 11693
rect 11498 11569 11601 11596
rect 11653 11569 11725 11596
rect 11777 11569 11849 11621
rect 11901 11569 11987 11621
rect 11498 11543 11987 11569
rect 393 10972 410 11543
rect 998 11125 1160 11136
rect 998 11079 1009 11125
rect 1149 11079 1160 11125
rect 998 11068 1160 11079
rect 2384 11125 2546 11136
rect 2384 11079 2395 11125
rect 2535 11079 2546 11125
rect 2384 11068 2546 11079
rect 2770 11125 2932 11136
rect 2770 11079 2781 11125
rect 2921 11079 2932 11125
rect 2770 11068 2932 11079
rect 4144 11125 4306 11136
rect 4144 11079 4155 11125
rect 4295 11079 4306 11125
rect 4144 11068 4306 11079
rect 4535 11125 4697 11136
rect 4535 11079 4546 11125
rect 4686 11079 4697 11125
rect 4535 11068 4697 11079
rect 5916 11125 6078 11136
rect 5916 11079 5927 11125
rect 6067 11079 6078 11125
rect 5916 11068 6078 11079
rect 6304 11125 6466 11136
rect 6304 11079 6315 11125
rect 6455 11079 6466 11125
rect 6304 11068 6466 11079
rect 7686 11125 7848 11136
rect 7686 11079 7697 11125
rect 7837 11079 7848 11125
rect 7686 11068 7848 11079
rect 8073 11125 8235 11136
rect 8073 11079 8084 11125
rect 8224 11079 8235 11125
rect 8073 11068 8235 11079
rect 9452 11125 9614 11136
rect 9452 11079 9463 11125
rect 9603 11079 9614 11125
rect 9452 11068 9614 11079
rect 9839 11125 10001 11136
rect 9839 11079 9850 11125
rect 9990 11079 10001 11125
rect 9839 11068 10001 11079
rect 11225 11125 11387 11136
rect 11225 11079 11236 11125
rect 11376 11079 11387 11125
rect 11225 11068 11387 11079
rect 393 10861 765 10972
rect 393 10289 440 10861
rect 700 10289 765 10861
rect 393 9852 765 10289
rect 393 7096 440 9852
rect 700 7096 765 9852
rect 393 6682 765 7096
rect 393 3926 440 6682
rect 700 3926 765 6682
rect 393 3505 765 3926
rect 393 3037 440 3505
rect 700 3037 765 3505
rect 393 2972 765 3037
rect 393 2420 410 2972
rect 1055 2876 1101 11068
rect 2441 2876 2487 11068
rect 2823 2876 2869 11068
rect 4209 2876 4255 11068
rect 4591 2876 4637 11068
rect 5977 2876 6023 11068
rect 6359 2876 6405 11068
rect 7745 2876 7791 11068
rect 8127 2876 8173 11068
rect 9513 2876 9559 11068
rect 9895 2876 9941 11068
rect 11281 2876 11327 11068
rect 11970 10972 11987 11543
rect 11615 10861 11987 10972
rect 11615 10289 11682 10861
rect 11942 10289 11987 10861
rect 11615 9852 11987 10289
rect 11615 7096 11682 9852
rect 11942 7096 11987 9852
rect 11615 6682 11987 7096
rect 11615 3926 11682 6682
rect 11942 3926 11987 6682
rect 11615 3505 11987 3926
rect 11615 3037 11682 3505
rect 11942 3037 11987 3505
rect 11615 2972 11987 3037
rect 998 2865 1160 2876
rect 998 2819 1009 2865
rect 1149 2819 1160 2865
rect 998 2808 1160 2819
rect 2384 2865 2546 2876
rect 2384 2819 2395 2865
rect 2535 2819 2546 2865
rect 2384 2808 2546 2819
rect 2770 2865 2932 2876
rect 2770 2819 2781 2865
rect 2921 2819 2932 2865
rect 2770 2808 2932 2819
rect 4144 2865 4306 2876
rect 4144 2819 4155 2865
rect 4295 2819 4306 2865
rect 4144 2808 4306 2819
rect 4535 2865 4697 2876
rect 4535 2819 4546 2865
rect 4686 2819 4697 2865
rect 4535 2808 4697 2819
rect 5916 2865 6078 2876
rect 5916 2819 5927 2865
rect 6067 2819 6078 2865
rect 5916 2808 6078 2819
rect 6304 2865 6466 2876
rect 6304 2819 6315 2865
rect 6455 2819 6466 2865
rect 6304 2808 6466 2819
rect 7686 2865 7848 2876
rect 7686 2819 7697 2865
rect 7837 2819 7848 2865
rect 7686 2808 7848 2819
rect 8073 2865 8235 2876
rect 8073 2819 8084 2865
rect 8224 2819 8235 2865
rect 8073 2808 8235 2819
rect 9452 2865 9614 2876
rect 9452 2819 9463 2865
rect 9603 2819 9614 2865
rect 9452 2808 9614 2819
rect 9839 2865 10001 2876
rect 9839 2819 9850 2865
rect 9990 2819 10001 2865
rect 9839 2808 10001 2819
rect 11225 2865 11387 2876
rect 11225 2819 11236 2865
rect 11376 2819 11387 2865
rect 11225 2808 11387 2819
rect 11970 2420 11987 2972
rect 393 2409 11987 2420
rect 393 2402 636 2409
rect 11782 2402 11987 2409
rect 393 2350 472 2402
rect 524 2350 596 2402
rect 11782 2350 11849 2402
rect 11901 2350 11987 2402
rect 393 2278 636 2350
rect 11782 2278 11987 2350
rect 393 2226 472 2278
rect 524 2226 596 2278
rect 11782 2226 11849 2278
rect 11901 2226 11987 2278
rect 393 2154 636 2226
rect 11782 2154 11987 2226
rect 393 2102 472 2154
rect 524 2102 596 2154
rect 11782 2102 11849 2154
rect 11901 2102 11987 2154
rect 393 2030 636 2102
rect 11782 2030 11987 2102
rect 393 1978 472 2030
rect 524 1978 596 2030
rect 11782 1978 11849 2030
rect 11901 1978 11987 2030
rect 393 1906 636 1978
rect 11782 1906 11987 1978
rect 393 1854 472 1906
rect 524 1854 596 1906
rect 11782 1854 11849 1906
rect 11901 1854 11987 1906
rect 393 1782 636 1854
rect 11782 1782 11987 1854
rect 393 1730 472 1782
rect 524 1730 596 1782
rect 11782 1730 11849 1782
rect 11901 1730 11987 1782
rect 393 1658 636 1730
rect 11782 1658 11987 1730
rect 393 1606 472 1658
rect 524 1606 596 1658
rect 11782 1606 11849 1658
rect 11901 1606 11987 1658
rect 393 1534 636 1606
rect 11782 1534 11987 1606
rect 393 1482 472 1534
rect 524 1482 596 1534
rect 11782 1482 11849 1534
rect 11901 1482 11987 1534
rect 393 1410 636 1482
rect 11782 1410 11987 1482
rect 393 1358 472 1410
rect 524 1358 596 1410
rect 11782 1358 11849 1410
rect 11901 1358 11987 1410
rect 393 1286 636 1358
rect 11782 1286 11987 1358
rect 393 1234 472 1286
rect 524 1234 596 1286
rect 11782 1234 11849 1286
rect 11901 1234 11987 1286
rect 393 1163 636 1234
rect 11782 1163 11987 1234
rect 393 1162 11987 1163
rect 393 1110 472 1162
rect 524 1110 596 1162
rect 648 1110 720 1162
rect 772 1110 11601 1162
rect 11653 1110 11725 1162
rect 11777 1110 11849 1162
rect 11901 1110 11987 1162
rect 393 1100 11987 1110
rect 12221 1100 12238 12990
rect 142 1061 12238 1100
rect 92 1038 12288 1061
rect 92 1014 472 1038
rect 524 1014 596 1038
rect 648 1014 720 1038
rect 772 1014 11601 1038
rect 11653 1014 11725 1038
rect 11777 1014 11849 1038
rect 11901 1014 12288 1038
rect 92 268 118 1014
rect 12264 268 12288 1014
rect 92 257 12288 268
rect 12444 52 12467 14481
rect -87 41 12467 52
rect -87 -805 118 41
rect 12264 -805 12467 41
rect -87 -865 12467 -805
rect 13113 -865 13136 14481
rect -756 -906 -696 -865
rect -540 -906 12891 -865
rect -756 -938 12891 -906
rect 13047 -938 13136 -865
rect -756 -1284 -733 -938
rect 13113 -1284 13136 -938
rect -756 -1301 13136 -1284
<< via1 >>
rect 466 15131 518 15183
rect 590 15131 642 15183
rect 714 15131 766 15183
rect 466 15007 518 15059
rect 590 15007 642 15059
rect 714 15007 766 15059
rect 466 14883 518 14935
rect 590 14883 642 14935
rect 714 14883 766 14935
rect 466 14759 518 14811
rect 590 14759 642 14811
rect 714 14759 766 14811
rect -719 14656 -667 14708
rect -611 14656 -559 14708
rect -503 14656 -451 14708
rect 466 14635 518 14687
rect 590 14635 642 14687
rect 714 14635 766 14687
rect -719 14593 -667 14600
rect -611 14593 -559 14600
rect -503 14593 -451 14600
rect -719 14548 -667 14593
rect -611 14548 -559 14593
rect -503 14548 -451 14593
rect -719 14481 -667 14492
rect -611 14481 -559 14492
rect -503 14481 -451 14492
rect -719 14440 -667 14481
rect -611 14440 -559 14481
rect -503 14440 -451 14481
rect -719 14332 -667 14384
rect -611 14332 -559 14384
rect -503 14332 -451 14384
rect -719 14224 -667 14276
rect -611 14224 -559 14276
rect -503 14224 -451 14276
rect -719 14116 -667 14168
rect -611 14116 -559 14168
rect -503 14116 -451 14168
rect -719 14008 -667 14060
rect -611 14008 -559 14060
rect -503 14008 -451 14060
rect -719 13900 -667 13952
rect -611 13900 -559 13952
rect -503 13900 -451 13952
rect -719 13792 -667 13844
rect -611 13792 -559 13844
rect -503 13792 -451 13844
rect -719 13684 -667 13736
rect -611 13684 -559 13736
rect -503 13684 -451 13736
rect -719 13576 -667 13628
rect -611 13576 -559 13628
rect -503 13576 -451 13628
rect -719 13468 -667 13520
rect -611 13468 -559 13520
rect -503 13468 -451 13520
rect -696 -865 -540 290
rect 1316 15147 1368 15199
rect 1440 15147 1492 15199
rect 1564 15147 1616 15199
rect 1688 15147 1740 15199
rect 1812 15147 1864 15199
rect 1936 15147 1988 15199
rect 2060 15147 2112 15199
rect 2184 15147 2236 15199
rect 1316 15023 1368 15075
rect 1440 15023 1492 15075
rect 1564 15023 1616 15075
rect 1688 15023 1740 15075
rect 1812 15023 1864 15075
rect 1936 15023 1988 15075
rect 2060 15023 2112 15075
rect 2184 15023 2236 15075
rect 1316 14899 1368 14951
rect 1440 14899 1492 14951
rect 1564 14899 1616 14951
rect 1688 14899 1740 14951
rect 1812 14899 1864 14951
rect 1936 14899 1988 14951
rect 2060 14899 2112 14951
rect 2184 14899 2236 14951
rect 1316 14775 1368 14827
rect 1440 14775 1492 14827
rect 1564 14775 1616 14827
rect 1688 14775 1740 14827
rect 1812 14775 1864 14827
rect 1936 14775 1988 14827
rect 2060 14775 2112 14827
rect 2184 14775 2236 14827
rect 1316 14651 1368 14703
rect 1440 14651 1492 14703
rect 1564 14651 1616 14703
rect 1688 14651 1740 14703
rect 1812 14651 1864 14703
rect 1936 14651 1988 14703
rect 2060 14651 2112 14703
rect 2184 14651 2236 14703
rect 1316 14527 1368 14579
rect 1440 14527 1492 14579
rect 1564 14527 1616 14579
rect 1688 14527 1740 14579
rect 1812 14527 1864 14579
rect 1936 14527 1988 14579
rect 2060 14527 2112 14579
rect 2184 14527 2236 14579
rect 1316 14403 1368 14455
rect 1440 14403 1492 14455
rect 1564 14403 1616 14455
rect 1688 14403 1740 14455
rect 1812 14403 1864 14455
rect 1936 14403 1988 14455
rect 2060 14403 2112 14455
rect 2184 14403 2236 14455
rect 3088 15147 3140 15199
rect 3212 15147 3264 15199
rect 3336 15147 3388 15199
rect 3460 15147 3512 15199
rect 3584 15147 3636 15199
rect 3708 15147 3760 15199
rect 3832 15147 3884 15199
rect 3956 15147 4008 15199
rect 3088 15023 3140 15075
rect 3212 15023 3264 15075
rect 3336 15023 3388 15075
rect 3460 15023 3512 15075
rect 3584 15023 3636 15075
rect 3708 15023 3760 15075
rect 3832 15023 3884 15075
rect 3956 15023 4008 15075
rect 3088 14899 3140 14951
rect 3212 14899 3264 14951
rect 3336 14899 3388 14951
rect 3460 14899 3512 14951
rect 3584 14899 3636 14951
rect 3708 14899 3760 14951
rect 3832 14899 3884 14951
rect 3956 14899 4008 14951
rect 3088 14775 3140 14827
rect 3212 14775 3264 14827
rect 3336 14775 3388 14827
rect 3460 14775 3512 14827
rect 3584 14775 3636 14827
rect 3708 14775 3760 14827
rect 3832 14775 3884 14827
rect 3956 14775 4008 14827
rect 3088 14651 3140 14703
rect 3212 14651 3264 14703
rect 3336 14651 3388 14703
rect 3460 14651 3512 14703
rect 3584 14651 3636 14703
rect 3708 14651 3760 14703
rect 3832 14651 3884 14703
rect 3956 14651 4008 14703
rect 3088 14527 3140 14579
rect 3212 14527 3264 14579
rect 3336 14527 3388 14579
rect 3460 14527 3512 14579
rect 3584 14527 3636 14579
rect 3708 14527 3760 14579
rect 3832 14527 3884 14579
rect 3956 14527 4008 14579
rect 3088 14403 3140 14455
rect 3212 14403 3264 14455
rect 3336 14403 3388 14455
rect 3460 14403 3512 14455
rect 3584 14403 3636 14455
rect 3708 14403 3760 14455
rect 3832 14403 3884 14455
rect 3956 14403 4008 14455
rect 4853 15147 4905 15199
rect 4977 15147 5029 15199
rect 5101 15147 5153 15199
rect 5225 15147 5277 15199
rect 5349 15147 5401 15199
rect 5473 15147 5525 15199
rect 5597 15147 5649 15199
rect 5721 15147 5773 15199
rect 4853 15023 4905 15075
rect 4977 15023 5029 15075
rect 5101 15023 5153 15075
rect 5225 15023 5277 15075
rect 5349 15023 5401 15075
rect 5473 15023 5525 15075
rect 5597 15023 5649 15075
rect 5721 15023 5773 15075
rect 4853 14899 4905 14951
rect 4977 14899 5029 14951
rect 5101 14899 5153 14951
rect 5225 14899 5277 14951
rect 5349 14899 5401 14951
rect 5473 14899 5525 14951
rect 5597 14899 5649 14951
rect 5721 14899 5773 14951
rect 4853 14775 4905 14827
rect 4977 14775 5029 14827
rect 5101 14775 5153 14827
rect 5225 14775 5277 14827
rect 5349 14775 5401 14827
rect 5473 14775 5525 14827
rect 5597 14775 5649 14827
rect 5721 14775 5773 14827
rect 4853 14651 4905 14703
rect 4977 14651 5029 14703
rect 5101 14651 5153 14703
rect 5225 14651 5277 14703
rect 5349 14651 5401 14703
rect 5473 14651 5525 14703
rect 5597 14651 5649 14703
rect 5721 14651 5773 14703
rect 4853 14527 4905 14579
rect 4977 14527 5029 14579
rect 5101 14527 5153 14579
rect 5225 14527 5277 14579
rect 5349 14527 5401 14579
rect 5473 14527 5525 14579
rect 5597 14527 5649 14579
rect 5721 14527 5773 14579
rect 4853 14403 4905 14455
rect 4977 14403 5029 14455
rect 5101 14403 5153 14455
rect 5225 14403 5277 14455
rect 5349 14403 5401 14455
rect 5473 14403 5525 14455
rect 5597 14403 5649 14455
rect 5721 14403 5773 14455
rect 6622 15147 6674 15199
rect 6746 15147 6798 15199
rect 6870 15147 6922 15199
rect 6994 15147 7046 15199
rect 7118 15147 7170 15199
rect 7242 15147 7294 15199
rect 7366 15147 7418 15199
rect 7490 15147 7542 15199
rect 6622 15023 6674 15075
rect 6746 15023 6798 15075
rect 6870 15023 6922 15075
rect 6994 15023 7046 15075
rect 7118 15023 7170 15075
rect 7242 15023 7294 15075
rect 7366 15023 7418 15075
rect 7490 15023 7542 15075
rect 6622 14899 6674 14951
rect 6746 14899 6798 14951
rect 6870 14899 6922 14951
rect 6994 14899 7046 14951
rect 7118 14899 7170 14951
rect 7242 14899 7294 14951
rect 7366 14899 7418 14951
rect 7490 14899 7542 14951
rect 6622 14775 6674 14827
rect 6746 14775 6798 14827
rect 6870 14775 6922 14827
rect 6994 14775 7046 14827
rect 7118 14775 7170 14827
rect 7242 14775 7294 14827
rect 7366 14775 7418 14827
rect 7490 14775 7542 14827
rect 6622 14651 6674 14703
rect 6746 14651 6798 14703
rect 6870 14651 6922 14703
rect 6994 14651 7046 14703
rect 7118 14651 7170 14703
rect 7242 14651 7294 14703
rect 7366 14651 7418 14703
rect 7490 14651 7542 14703
rect 6622 14527 6674 14579
rect 6746 14527 6798 14579
rect 6870 14527 6922 14579
rect 6994 14527 7046 14579
rect 7118 14527 7170 14579
rect 7242 14527 7294 14579
rect 7366 14527 7418 14579
rect 7490 14527 7542 14579
rect 6622 14403 6674 14455
rect 6746 14403 6798 14455
rect 6870 14403 6922 14455
rect 6994 14403 7046 14455
rect 7118 14403 7170 14455
rect 7242 14403 7294 14455
rect 7366 14403 7418 14455
rect 7490 14403 7542 14455
rect 8391 15147 8443 15199
rect 8515 15147 8567 15199
rect 8639 15147 8691 15199
rect 8763 15147 8815 15199
rect 8887 15147 8939 15199
rect 9011 15147 9063 15199
rect 9135 15147 9187 15199
rect 9259 15147 9311 15199
rect 8391 15023 8443 15075
rect 8515 15023 8567 15075
rect 8639 15023 8691 15075
rect 8763 15023 8815 15075
rect 8887 15023 8939 15075
rect 9011 15023 9063 15075
rect 9135 15023 9187 15075
rect 9259 15023 9311 15075
rect 8391 14899 8443 14951
rect 8515 14899 8567 14951
rect 8639 14899 8691 14951
rect 8763 14899 8815 14951
rect 8887 14899 8939 14951
rect 9011 14899 9063 14951
rect 9135 14899 9187 14951
rect 9259 14899 9311 14951
rect 8391 14775 8443 14827
rect 8515 14775 8567 14827
rect 8639 14775 8691 14827
rect 8763 14775 8815 14827
rect 8887 14775 8939 14827
rect 9011 14775 9063 14827
rect 9135 14775 9187 14827
rect 9259 14775 9311 14827
rect 8391 14651 8443 14703
rect 8515 14651 8567 14703
rect 8639 14651 8691 14703
rect 8763 14651 8815 14703
rect 8887 14651 8939 14703
rect 9011 14651 9063 14703
rect 9135 14651 9187 14703
rect 9259 14651 9311 14703
rect 8391 14527 8443 14579
rect 8515 14527 8567 14579
rect 8639 14527 8691 14579
rect 8763 14527 8815 14579
rect 8887 14527 8939 14579
rect 9011 14527 9063 14579
rect 9135 14527 9187 14579
rect 9259 14527 9311 14579
rect 8391 14403 8443 14455
rect 8515 14403 8567 14455
rect 8639 14403 8691 14455
rect 8763 14403 8815 14455
rect 8887 14403 8939 14455
rect 9011 14403 9063 14455
rect 9135 14403 9187 14455
rect 9259 14403 9311 14455
rect 10157 15147 10209 15199
rect 10281 15147 10333 15199
rect 10405 15147 10457 15199
rect 10529 15147 10581 15199
rect 10653 15147 10705 15199
rect 10777 15147 10829 15199
rect 10901 15147 10953 15199
rect 11025 15147 11077 15199
rect 10157 15023 10209 15075
rect 10281 15023 10333 15075
rect 10405 15023 10457 15075
rect 10529 15023 10581 15075
rect 10653 15023 10705 15075
rect 10777 15023 10829 15075
rect 10901 15023 10953 15075
rect 11025 15023 11077 15075
rect 10157 14899 10209 14951
rect 10281 14899 10333 14951
rect 10405 14899 10457 14951
rect 10529 14899 10581 14951
rect 10653 14899 10705 14951
rect 10777 14899 10829 14951
rect 10901 14899 10953 14951
rect 11025 14899 11077 14951
rect 10157 14775 10209 14827
rect 10281 14775 10333 14827
rect 10405 14775 10457 14827
rect 10529 14775 10581 14827
rect 10653 14775 10705 14827
rect 10777 14775 10829 14827
rect 10901 14775 10953 14827
rect 11025 14775 11077 14827
rect 10157 14651 10209 14703
rect 10281 14651 10333 14703
rect 10405 14651 10457 14703
rect 10529 14651 10581 14703
rect 10653 14651 10705 14703
rect 10777 14651 10829 14703
rect 10901 14651 10953 14703
rect 11025 14651 11077 14703
rect 10157 14527 10209 14579
rect 10281 14527 10333 14579
rect 10405 14527 10457 14579
rect 10529 14527 10581 14579
rect 10653 14527 10705 14579
rect 10777 14527 10829 14579
rect 10901 14527 10953 14579
rect 11025 14527 11077 14579
rect 10157 14403 10209 14455
rect 10281 14403 10333 14455
rect 10405 14403 10457 14455
rect 10529 14403 10581 14455
rect 10653 14403 10705 14455
rect 10777 14403 10829 14455
rect 10901 14403 10953 14455
rect 11025 14403 11077 14455
rect 11595 15131 11647 15183
rect 11719 15131 11771 15183
rect 11843 15131 11895 15183
rect 11595 15007 11647 15059
rect 11719 15007 11771 15059
rect 11843 15007 11895 15059
rect 11595 14883 11647 14935
rect 11719 14883 11771 14935
rect 11843 14883 11895 14935
rect 11595 14759 11647 14811
rect 11719 14759 11771 14811
rect 11843 14759 11895 14811
rect 11595 14635 11647 14687
rect 11719 14635 11771 14687
rect 11843 14635 11895 14687
rect 472 13057 524 13109
rect 596 13057 648 13109
rect 720 13057 772 13109
rect 472 12933 524 12985
rect 596 12958 648 12985
rect 720 12958 772 12985
rect 596 12933 624 12958
rect 624 12933 648 12958
rect 720 12933 772 12958
rect 472 12809 524 12861
rect 596 12809 624 12861
rect 624 12809 648 12861
rect 720 12809 772 12861
rect 472 12685 524 12737
rect 596 12685 624 12737
rect 624 12685 648 12737
rect 720 12685 772 12737
rect 472 12561 524 12613
rect 596 12561 624 12613
rect 624 12561 648 12613
rect 720 12561 772 12613
rect 472 12437 524 12489
rect 596 12437 624 12489
rect 624 12437 648 12489
rect 720 12437 772 12489
rect 472 12313 524 12365
rect 596 12313 624 12365
rect 624 12313 648 12365
rect 720 12313 772 12365
rect 472 12189 524 12241
rect 596 12189 624 12241
rect 624 12189 648 12241
rect 720 12189 772 12241
rect 472 12065 524 12117
rect 596 12065 624 12117
rect 624 12065 648 12117
rect 720 12065 772 12117
rect 472 11941 524 11993
rect 596 11941 624 11993
rect 624 11941 648 11993
rect 720 11941 772 11993
rect 472 11817 524 11869
rect 596 11817 624 11869
rect 624 11817 648 11869
rect 720 11817 772 11869
rect 472 11693 524 11745
rect 596 11693 624 11745
rect 624 11693 648 11745
rect 720 11693 772 11745
rect 472 11569 524 11621
rect 596 11596 624 11621
rect 624 11596 648 11621
rect 720 11596 772 11621
rect 596 11569 648 11596
rect 720 11569 772 11596
rect 11601 13057 11653 13109
rect 11725 13057 11777 13109
rect 11849 13057 11901 13109
rect 11601 12958 11653 12985
rect 11725 12958 11777 12985
rect 11601 12933 11653 12958
rect 11725 12933 11758 12958
rect 11758 12933 11777 12958
rect 11849 12933 11901 12985
rect 11601 12809 11653 12861
rect 11725 12809 11758 12861
rect 11758 12809 11777 12861
rect 11849 12809 11901 12861
rect 11601 12685 11653 12737
rect 11725 12685 11758 12737
rect 11758 12685 11777 12737
rect 11849 12685 11901 12737
rect 11601 12561 11653 12613
rect 11725 12561 11758 12613
rect 11758 12561 11777 12613
rect 11849 12561 11901 12613
rect 11601 12437 11653 12489
rect 11725 12437 11758 12489
rect 11758 12437 11777 12489
rect 11849 12437 11901 12489
rect 11601 12313 11653 12365
rect 11725 12313 11758 12365
rect 11758 12313 11777 12365
rect 11849 12313 11901 12365
rect 11601 12189 11653 12241
rect 11725 12189 11758 12241
rect 11758 12189 11777 12241
rect 11849 12189 11901 12241
rect 11601 12065 11653 12117
rect 11725 12065 11758 12117
rect 11758 12065 11777 12117
rect 11849 12065 11901 12117
rect 11601 11941 11653 11993
rect 11725 11941 11758 11993
rect 11758 11941 11777 11993
rect 11849 11941 11901 11993
rect 11601 11817 11653 11869
rect 11725 11817 11758 11869
rect 11758 11817 11777 11869
rect 11849 11817 11901 11869
rect 11601 11693 11653 11745
rect 11725 11693 11758 11745
rect 11758 11693 11777 11745
rect 11849 11693 11901 11745
rect 11601 11596 11653 11621
rect 11725 11596 11758 11621
rect 11758 11596 11777 11621
rect 11601 11569 11653 11596
rect 11725 11569 11777 11596
rect 11849 11569 11901 11621
rect 440 10289 700 10861
rect 440 7096 700 9852
rect 440 3926 700 6682
rect 440 3037 700 3505
rect 11682 10289 11942 10861
rect 11682 7096 11942 9852
rect 11682 3926 11942 6682
rect 11682 3037 11942 3505
rect 472 2350 524 2402
rect 596 2350 636 2402
rect 636 2350 648 2402
rect 720 2350 772 2402
rect 11601 2350 11653 2402
rect 11725 2350 11777 2402
rect 11849 2350 11901 2402
rect 472 2226 524 2278
rect 596 2226 636 2278
rect 636 2226 648 2278
rect 720 2226 772 2278
rect 11601 2226 11653 2278
rect 11725 2226 11777 2278
rect 11849 2226 11901 2278
rect 472 2102 524 2154
rect 596 2102 636 2154
rect 636 2102 648 2154
rect 720 2102 772 2154
rect 11601 2102 11653 2154
rect 11725 2102 11777 2154
rect 11849 2102 11901 2154
rect 472 1978 524 2030
rect 596 1978 636 2030
rect 636 1978 648 2030
rect 720 1978 772 2030
rect 11601 1978 11653 2030
rect 11725 1978 11777 2030
rect 11849 1978 11901 2030
rect 472 1854 524 1906
rect 596 1854 636 1906
rect 636 1854 648 1906
rect 720 1854 772 1906
rect 11601 1854 11653 1906
rect 11725 1854 11777 1906
rect 11849 1854 11901 1906
rect 472 1730 524 1782
rect 596 1730 636 1782
rect 636 1730 648 1782
rect 720 1730 772 1782
rect 11601 1730 11653 1782
rect 11725 1730 11777 1782
rect 11849 1730 11901 1782
rect 472 1606 524 1658
rect 596 1606 636 1658
rect 636 1606 648 1658
rect 720 1606 772 1658
rect 11601 1606 11653 1658
rect 11725 1606 11777 1658
rect 11849 1606 11901 1658
rect 472 1482 524 1534
rect 596 1482 636 1534
rect 636 1482 648 1534
rect 720 1482 772 1534
rect 11601 1482 11653 1534
rect 11725 1482 11777 1534
rect 11849 1482 11901 1534
rect 472 1358 524 1410
rect 596 1358 636 1410
rect 636 1358 648 1410
rect 720 1358 772 1410
rect 11601 1358 11653 1410
rect 11725 1358 11777 1410
rect 11849 1358 11901 1410
rect 472 1234 524 1286
rect 596 1234 636 1286
rect 636 1234 648 1286
rect 720 1234 772 1286
rect 11601 1234 11653 1286
rect 11725 1234 11777 1286
rect 11849 1234 11901 1286
rect 472 1110 524 1162
rect 596 1110 648 1162
rect 720 1110 772 1162
rect 11601 1110 11653 1162
rect 11725 1110 11777 1162
rect 11849 1110 11901 1162
rect 472 1014 524 1038
rect 596 1014 648 1038
rect 720 1014 772 1038
rect 11601 1014 11653 1038
rect 11725 1014 11777 1038
rect 11849 1014 11901 1038
rect 472 986 524 1014
rect 596 986 648 1014
rect 720 986 772 1014
rect 11601 986 11653 1014
rect 11725 986 11777 1014
rect 11849 986 11901 1014
rect 472 862 524 914
rect 596 862 648 914
rect 720 862 772 914
rect 11601 862 11653 914
rect 11725 862 11777 914
rect 11849 862 11901 914
rect 472 738 524 790
rect 596 738 648 790
rect 720 738 772 790
rect 11601 738 11653 790
rect 11725 738 11777 790
rect 11849 738 11901 790
rect 472 614 524 666
rect 596 614 648 666
rect 720 614 772 666
rect 11601 614 11653 666
rect 11725 614 11777 666
rect 11849 614 11901 666
rect 12891 -865 13047 339
rect -696 -906 -540 -865
rect 12891 -938 13047 -865
rect 12891 -961 13047 -938
<< metal2 >>
rect 416 15183 816 15250
rect 416 15131 466 15183
rect 518 15131 590 15183
rect 642 15131 714 15183
rect 766 15131 816 15183
rect 416 15059 816 15131
rect 416 15007 466 15059
rect 518 15007 590 15059
rect 642 15007 714 15059
rect 766 15007 816 15059
rect 416 14935 816 15007
rect 416 14883 466 14935
rect 518 14883 590 14935
rect 642 14883 714 14935
rect 766 14883 816 14935
rect -756 14755 -439 14820
rect -756 14708 -684 14755
rect -628 14708 -542 14755
rect -486 14708 -439 14755
rect -756 14656 -719 14708
rect -628 14699 -611 14708
rect -667 14656 -611 14699
rect -559 14699 -542 14708
rect -559 14656 -503 14699
rect -451 14656 -439 14708
rect -756 14613 -439 14656
rect -756 14600 -684 14613
rect -628 14600 -542 14613
rect -486 14600 -439 14613
rect -756 14548 -719 14600
rect -628 14557 -611 14600
rect -667 14548 -611 14557
rect -559 14557 -542 14600
rect -559 14548 -503 14557
rect -451 14548 -439 14600
rect -756 14492 -439 14548
rect -756 14440 -719 14492
rect -667 14471 -611 14492
rect -628 14440 -611 14471
rect -559 14471 -503 14492
rect -559 14440 -542 14471
rect -451 14440 -439 14492
rect -756 14415 -684 14440
rect -628 14415 -542 14440
rect -486 14415 -439 14440
rect -756 14384 -439 14415
rect -756 14332 -719 14384
rect -667 14332 -611 14384
rect -559 14332 -503 14384
rect -451 14332 -439 14384
rect -756 14329 -439 14332
rect -756 14276 -684 14329
rect -628 14276 -542 14329
rect -486 14276 -439 14329
rect -756 14224 -719 14276
rect -628 14273 -611 14276
rect -667 14224 -611 14273
rect -559 14273 -542 14276
rect -559 14224 -503 14273
rect -451 14224 -439 14276
rect -756 14187 -439 14224
rect -756 14168 -684 14187
rect -628 14168 -542 14187
rect -486 14168 -439 14187
rect -756 14116 -719 14168
rect -628 14131 -611 14168
rect -667 14116 -611 14131
rect -559 14131 -542 14168
rect -559 14116 -503 14131
rect -451 14116 -439 14168
rect -756 14060 -439 14116
rect -756 14008 -719 14060
rect -667 14045 -611 14060
rect -628 14008 -611 14045
rect -559 14045 -503 14060
rect -559 14008 -542 14045
rect -451 14008 -439 14060
rect -756 13989 -684 14008
rect -628 13989 -542 14008
rect -486 13989 -439 14008
rect -756 13952 -439 13989
rect -756 13900 -719 13952
rect -667 13903 -611 13952
rect -628 13900 -611 13903
rect -559 13903 -503 13952
rect -559 13900 -542 13903
rect -451 13900 -439 13952
rect -756 13847 -684 13900
rect -628 13847 -542 13900
rect -486 13847 -439 13900
rect -756 13844 -439 13847
rect -756 13792 -719 13844
rect -667 13792 -611 13844
rect -559 13792 -503 13844
rect -451 13792 -439 13844
rect -756 13761 -439 13792
rect -756 13736 -684 13761
rect -628 13736 -542 13761
rect -486 13736 -439 13761
rect -756 13684 -719 13736
rect -628 13705 -611 13736
rect -667 13684 -611 13705
rect -559 13705 -542 13736
rect -559 13684 -503 13705
rect -451 13684 -439 13736
rect -756 13628 -439 13684
rect -756 13576 -719 13628
rect -667 13619 -611 13628
rect -628 13576 -611 13619
rect -559 13619 -503 13628
rect -559 13576 -542 13619
rect -451 13576 -439 13628
rect -756 13563 -684 13576
rect -628 13563 -542 13576
rect -486 13563 -439 13576
rect -756 13520 -439 13563
rect -756 13468 -719 13520
rect -667 13477 -611 13520
rect -628 13468 -611 13477
rect -559 13477 -503 13520
rect -559 13468 -542 13477
rect -451 13468 -439 13520
rect -756 13421 -684 13468
rect -628 13421 -542 13468
rect -486 13421 -439 13468
rect -756 13411 -439 13421
rect 416 14811 816 14883
rect 416 14759 466 14811
rect 518 14759 590 14811
rect 642 14759 714 14811
rect 766 14759 816 14811
rect 416 14755 816 14759
rect 416 14699 446 14755
rect 502 14699 588 14755
rect 644 14699 730 14755
rect 786 14699 816 14755
rect 416 14687 816 14699
rect 416 14635 466 14687
rect 518 14635 590 14687
rect 642 14635 714 14687
rect 766 14635 816 14687
rect 416 14613 816 14635
rect 416 14557 446 14613
rect 502 14557 588 14613
rect 644 14557 730 14613
rect 786 14557 816 14613
rect 416 14471 816 14557
rect 416 14415 446 14471
rect 502 14415 588 14471
rect 644 14415 730 14471
rect 786 14415 816 14471
rect 416 14329 816 14415
rect 1304 15199 2248 15211
rect 1304 15147 1316 15199
rect 1368 15147 1440 15199
rect 1492 15147 1564 15199
rect 1616 15147 1688 15199
rect 1740 15147 1812 15199
rect 1864 15147 1936 15199
rect 1988 15147 2060 15199
rect 2112 15147 2184 15199
rect 2236 15147 2248 15199
rect 1304 15075 2248 15147
rect 1304 15023 1316 15075
rect 1368 15023 1440 15075
rect 1492 15023 1564 15075
rect 1616 15023 1688 15075
rect 1740 15023 1812 15075
rect 1864 15023 1936 15075
rect 1988 15023 2060 15075
rect 2112 15023 2184 15075
rect 2236 15023 2248 15075
rect 1304 14951 2248 15023
rect 1304 14899 1316 14951
rect 1368 14899 1440 14951
rect 1492 14899 1564 14951
rect 1616 14899 1688 14951
rect 1740 14899 1812 14951
rect 1864 14899 1936 14951
rect 1988 14899 2060 14951
rect 2112 14899 2184 14951
rect 2236 14899 2248 14951
rect 1304 14827 2248 14899
rect 1304 14775 1316 14827
rect 1368 14775 1440 14827
rect 1492 14775 1564 14827
rect 1616 14775 1688 14827
rect 1740 14775 1812 14827
rect 1864 14775 1936 14827
rect 1988 14775 2060 14827
rect 2112 14775 2184 14827
rect 2236 14775 2248 14827
rect 1304 14748 2248 14775
rect 1304 14703 1322 14748
rect 1378 14703 1464 14748
rect 1520 14703 1606 14748
rect 1662 14703 1748 14748
rect 1304 14651 1316 14703
rect 1378 14692 1440 14703
rect 1520 14692 1564 14703
rect 1662 14692 1688 14703
rect 1368 14651 1440 14692
rect 1492 14651 1564 14692
rect 1616 14651 1688 14692
rect 1740 14692 1748 14703
rect 1804 14703 1890 14748
rect 1946 14703 2032 14748
rect 2088 14703 2174 14748
rect 2230 14703 2248 14748
rect 1804 14692 1812 14703
rect 1740 14651 1812 14692
rect 1864 14692 1890 14703
rect 1988 14692 2032 14703
rect 2112 14692 2174 14703
rect 1864 14651 1936 14692
rect 1988 14651 2060 14692
rect 2112 14651 2184 14692
rect 2236 14651 2248 14703
rect 1304 14606 2248 14651
rect 1304 14579 1322 14606
rect 1378 14579 1464 14606
rect 1520 14579 1606 14606
rect 1662 14579 1748 14606
rect 1304 14527 1316 14579
rect 1378 14550 1440 14579
rect 1520 14550 1564 14579
rect 1662 14550 1688 14579
rect 1368 14527 1440 14550
rect 1492 14527 1564 14550
rect 1616 14527 1688 14550
rect 1740 14550 1748 14579
rect 1804 14579 1890 14606
rect 1946 14579 2032 14606
rect 2088 14579 2174 14606
rect 2230 14579 2248 14606
rect 1804 14550 1812 14579
rect 1740 14527 1812 14550
rect 1864 14550 1890 14579
rect 1988 14550 2032 14579
rect 2112 14550 2174 14579
rect 1864 14527 1936 14550
rect 1988 14527 2060 14550
rect 2112 14527 2184 14550
rect 2236 14527 2248 14579
rect 1304 14464 2248 14527
rect 1304 14455 1322 14464
rect 1378 14455 1464 14464
rect 1520 14455 1606 14464
rect 1662 14455 1748 14464
rect 1304 14403 1316 14455
rect 1378 14408 1440 14455
rect 1520 14408 1564 14455
rect 1662 14408 1688 14455
rect 1368 14403 1440 14408
rect 1492 14403 1564 14408
rect 1616 14403 1688 14408
rect 1740 14408 1748 14455
rect 1804 14455 1890 14464
rect 1946 14455 2032 14464
rect 2088 14455 2174 14464
rect 2230 14455 2248 14464
rect 1804 14408 1812 14455
rect 1740 14403 1812 14408
rect 1864 14408 1890 14455
rect 1988 14408 2032 14455
rect 2112 14408 2174 14455
rect 1864 14403 1936 14408
rect 1988 14403 2060 14408
rect 2112 14403 2184 14408
rect 2236 14403 2248 14455
rect 1304 14391 2248 14403
rect 3076 15199 4020 15211
rect 3076 15147 3088 15199
rect 3140 15147 3212 15199
rect 3264 15147 3336 15199
rect 3388 15147 3460 15199
rect 3512 15147 3584 15199
rect 3636 15147 3708 15199
rect 3760 15147 3832 15199
rect 3884 15147 3956 15199
rect 4008 15147 4020 15199
rect 3076 15075 4020 15147
rect 3076 15023 3088 15075
rect 3140 15023 3212 15075
rect 3264 15023 3336 15075
rect 3388 15023 3460 15075
rect 3512 15023 3584 15075
rect 3636 15023 3708 15075
rect 3760 15023 3832 15075
rect 3884 15023 3956 15075
rect 4008 15023 4020 15075
rect 3076 14951 4020 15023
rect 3076 14899 3088 14951
rect 3140 14899 3212 14951
rect 3264 14899 3336 14951
rect 3388 14899 3460 14951
rect 3512 14899 3584 14951
rect 3636 14899 3708 14951
rect 3760 14899 3832 14951
rect 3884 14899 3956 14951
rect 4008 14899 4020 14951
rect 3076 14827 4020 14899
rect 3076 14775 3088 14827
rect 3140 14775 3212 14827
rect 3264 14775 3336 14827
rect 3388 14775 3460 14827
rect 3512 14775 3584 14827
rect 3636 14775 3708 14827
rect 3760 14775 3832 14827
rect 3884 14775 3956 14827
rect 4008 14775 4020 14827
rect 3076 14748 4020 14775
rect 3076 14703 3094 14748
rect 3150 14703 3236 14748
rect 3292 14703 3378 14748
rect 3434 14703 3520 14748
rect 3076 14651 3088 14703
rect 3150 14692 3212 14703
rect 3292 14692 3336 14703
rect 3434 14692 3460 14703
rect 3140 14651 3212 14692
rect 3264 14651 3336 14692
rect 3388 14651 3460 14692
rect 3512 14692 3520 14703
rect 3576 14703 3662 14748
rect 3718 14703 3804 14748
rect 3860 14703 3946 14748
rect 4002 14703 4020 14748
rect 3576 14692 3584 14703
rect 3512 14651 3584 14692
rect 3636 14692 3662 14703
rect 3760 14692 3804 14703
rect 3884 14692 3946 14703
rect 3636 14651 3708 14692
rect 3760 14651 3832 14692
rect 3884 14651 3956 14692
rect 4008 14651 4020 14703
rect 3076 14606 4020 14651
rect 3076 14579 3094 14606
rect 3150 14579 3236 14606
rect 3292 14579 3378 14606
rect 3434 14579 3520 14606
rect 3076 14527 3088 14579
rect 3150 14550 3212 14579
rect 3292 14550 3336 14579
rect 3434 14550 3460 14579
rect 3140 14527 3212 14550
rect 3264 14527 3336 14550
rect 3388 14527 3460 14550
rect 3512 14550 3520 14579
rect 3576 14579 3662 14606
rect 3718 14579 3804 14606
rect 3860 14579 3946 14606
rect 4002 14579 4020 14606
rect 3576 14550 3584 14579
rect 3512 14527 3584 14550
rect 3636 14550 3662 14579
rect 3760 14550 3804 14579
rect 3884 14550 3946 14579
rect 3636 14527 3708 14550
rect 3760 14527 3832 14550
rect 3884 14527 3956 14550
rect 4008 14527 4020 14579
rect 3076 14464 4020 14527
rect 3076 14455 3094 14464
rect 3150 14455 3236 14464
rect 3292 14455 3378 14464
rect 3434 14455 3520 14464
rect 3076 14403 3088 14455
rect 3150 14408 3212 14455
rect 3292 14408 3336 14455
rect 3434 14408 3460 14455
rect 3140 14403 3212 14408
rect 3264 14403 3336 14408
rect 3388 14403 3460 14408
rect 3512 14408 3520 14455
rect 3576 14455 3662 14464
rect 3718 14455 3804 14464
rect 3860 14455 3946 14464
rect 4002 14455 4020 14464
rect 3576 14408 3584 14455
rect 3512 14403 3584 14408
rect 3636 14408 3662 14455
rect 3760 14408 3804 14455
rect 3884 14408 3946 14455
rect 3636 14403 3708 14408
rect 3760 14403 3832 14408
rect 3884 14403 3956 14408
rect 4008 14403 4020 14455
rect 3076 14391 4020 14403
rect 4841 15199 5785 15211
rect 4841 15147 4853 15199
rect 4905 15147 4977 15199
rect 5029 15147 5101 15199
rect 5153 15147 5225 15199
rect 5277 15147 5349 15199
rect 5401 15147 5473 15199
rect 5525 15147 5597 15199
rect 5649 15147 5721 15199
rect 5773 15147 5785 15199
rect 4841 15075 5785 15147
rect 4841 15023 4853 15075
rect 4905 15023 4977 15075
rect 5029 15023 5101 15075
rect 5153 15023 5225 15075
rect 5277 15023 5349 15075
rect 5401 15023 5473 15075
rect 5525 15023 5597 15075
rect 5649 15023 5721 15075
rect 5773 15023 5785 15075
rect 4841 14951 5785 15023
rect 4841 14899 4853 14951
rect 4905 14899 4977 14951
rect 5029 14899 5101 14951
rect 5153 14899 5225 14951
rect 5277 14899 5349 14951
rect 5401 14899 5473 14951
rect 5525 14899 5597 14951
rect 5649 14899 5721 14951
rect 5773 14899 5785 14951
rect 4841 14827 5785 14899
rect 4841 14775 4853 14827
rect 4905 14775 4977 14827
rect 5029 14775 5101 14827
rect 5153 14775 5225 14827
rect 5277 14775 5349 14827
rect 5401 14775 5473 14827
rect 5525 14775 5597 14827
rect 5649 14775 5721 14827
rect 5773 14775 5785 14827
rect 4841 14748 5785 14775
rect 4841 14703 4859 14748
rect 4915 14703 5001 14748
rect 5057 14703 5143 14748
rect 5199 14703 5285 14748
rect 4841 14651 4853 14703
rect 4915 14692 4977 14703
rect 5057 14692 5101 14703
rect 5199 14692 5225 14703
rect 4905 14651 4977 14692
rect 5029 14651 5101 14692
rect 5153 14651 5225 14692
rect 5277 14692 5285 14703
rect 5341 14703 5427 14748
rect 5483 14703 5569 14748
rect 5625 14703 5711 14748
rect 5767 14703 5785 14748
rect 5341 14692 5349 14703
rect 5277 14651 5349 14692
rect 5401 14692 5427 14703
rect 5525 14692 5569 14703
rect 5649 14692 5711 14703
rect 5401 14651 5473 14692
rect 5525 14651 5597 14692
rect 5649 14651 5721 14692
rect 5773 14651 5785 14703
rect 4841 14606 5785 14651
rect 4841 14579 4859 14606
rect 4915 14579 5001 14606
rect 5057 14579 5143 14606
rect 5199 14579 5285 14606
rect 4841 14527 4853 14579
rect 4915 14550 4977 14579
rect 5057 14550 5101 14579
rect 5199 14550 5225 14579
rect 4905 14527 4977 14550
rect 5029 14527 5101 14550
rect 5153 14527 5225 14550
rect 5277 14550 5285 14579
rect 5341 14579 5427 14606
rect 5483 14579 5569 14606
rect 5625 14579 5711 14606
rect 5767 14579 5785 14606
rect 5341 14550 5349 14579
rect 5277 14527 5349 14550
rect 5401 14550 5427 14579
rect 5525 14550 5569 14579
rect 5649 14550 5711 14579
rect 5401 14527 5473 14550
rect 5525 14527 5597 14550
rect 5649 14527 5721 14550
rect 5773 14527 5785 14579
rect 4841 14464 5785 14527
rect 4841 14455 4859 14464
rect 4915 14455 5001 14464
rect 5057 14455 5143 14464
rect 5199 14455 5285 14464
rect 4841 14403 4853 14455
rect 4915 14408 4977 14455
rect 5057 14408 5101 14455
rect 5199 14408 5225 14455
rect 4905 14403 4977 14408
rect 5029 14403 5101 14408
rect 5153 14403 5225 14408
rect 5277 14408 5285 14455
rect 5341 14455 5427 14464
rect 5483 14455 5569 14464
rect 5625 14455 5711 14464
rect 5767 14455 5785 14464
rect 5341 14408 5349 14455
rect 5277 14403 5349 14408
rect 5401 14408 5427 14455
rect 5525 14408 5569 14455
rect 5649 14408 5711 14455
rect 5401 14403 5473 14408
rect 5525 14403 5597 14408
rect 5649 14403 5721 14408
rect 5773 14403 5785 14455
rect 4841 14391 5785 14403
rect 6610 15199 7554 15211
rect 6610 15147 6622 15199
rect 6674 15147 6746 15199
rect 6798 15147 6870 15199
rect 6922 15147 6994 15199
rect 7046 15147 7118 15199
rect 7170 15147 7242 15199
rect 7294 15147 7366 15199
rect 7418 15147 7490 15199
rect 7542 15147 7554 15199
rect 6610 15075 7554 15147
rect 6610 15023 6622 15075
rect 6674 15023 6746 15075
rect 6798 15023 6870 15075
rect 6922 15023 6994 15075
rect 7046 15023 7118 15075
rect 7170 15023 7242 15075
rect 7294 15023 7366 15075
rect 7418 15023 7490 15075
rect 7542 15023 7554 15075
rect 6610 14951 7554 15023
rect 6610 14899 6622 14951
rect 6674 14899 6746 14951
rect 6798 14899 6870 14951
rect 6922 14899 6994 14951
rect 7046 14899 7118 14951
rect 7170 14899 7242 14951
rect 7294 14899 7366 14951
rect 7418 14899 7490 14951
rect 7542 14899 7554 14951
rect 6610 14827 7554 14899
rect 6610 14775 6622 14827
rect 6674 14775 6746 14827
rect 6798 14775 6870 14827
rect 6922 14775 6994 14827
rect 7046 14775 7118 14827
rect 7170 14775 7242 14827
rect 7294 14775 7366 14827
rect 7418 14775 7490 14827
rect 7542 14775 7554 14827
rect 6610 14748 7554 14775
rect 6610 14703 6628 14748
rect 6684 14703 6770 14748
rect 6826 14703 6912 14748
rect 6968 14703 7054 14748
rect 6610 14651 6622 14703
rect 6684 14692 6746 14703
rect 6826 14692 6870 14703
rect 6968 14692 6994 14703
rect 6674 14651 6746 14692
rect 6798 14651 6870 14692
rect 6922 14651 6994 14692
rect 7046 14692 7054 14703
rect 7110 14703 7196 14748
rect 7252 14703 7338 14748
rect 7394 14703 7480 14748
rect 7536 14703 7554 14748
rect 7110 14692 7118 14703
rect 7046 14651 7118 14692
rect 7170 14692 7196 14703
rect 7294 14692 7338 14703
rect 7418 14692 7480 14703
rect 7170 14651 7242 14692
rect 7294 14651 7366 14692
rect 7418 14651 7490 14692
rect 7542 14651 7554 14703
rect 6610 14606 7554 14651
rect 6610 14579 6628 14606
rect 6684 14579 6770 14606
rect 6826 14579 6912 14606
rect 6968 14579 7054 14606
rect 6610 14527 6622 14579
rect 6684 14550 6746 14579
rect 6826 14550 6870 14579
rect 6968 14550 6994 14579
rect 6674 14527 6746 14550
rect 6798 14527 6870 14550
rect 6922 14527 6994 14550
rect 7046 14550 7054 14579
rect 7110 14579 7196 14606
rect 7252 14579 7338 14606
rect 7394 14579 7480 14606
rect 7536 14579 7554 14606
rect 7110 14550 7118 14579
rect 7046 14527 7118 14550
rect 7170 14550 7196 14579
rect 7294 14550 7338 14579
rect 7418 14550 7480 14579
rect 7170 14527 7242 14550
rect 7294 14527 7366 14550
rect 7418 14527 7490 14550
rect 7542 14527 7554 14579
rect 6610 14464 7554 14527
rect 6610 14455 6628 14464
rect 6684 14455 6770 14464
rect 6826 14455 6912 14464
rect 6968 14455 7054 14464
rect 6610 14403 6622 14455
rect 6684 14408 6746 14455
rect 6826 14408 6870 14455
rect 6968 14408 6994 14455
rect 6674 14403 6746 14408
rect 6798 14403 6870 14408
rect 6922 14403 6994 14408
rect 7046 14408 7054 14455
rect 7110 14455 7196 14464
rect 7252 14455 7338 14464
rect 7394 14455 7480 14464
rect 7536 14455 7554 14464
rect 7110 14408 7118 14455
rect 7046 14403 7118 14408
rect 7170 14408 7196 14455
rect 7294 14408 7338 14455
rect 7418 14408 7480 14455
rect 7170 14403 7242 14408
rect 7294 14403 7366 14408
rect 7418 14403 7490 14408
rect 7542 14403 7554 14455
rect 6610 14391 7554 14403
rect 8379 15199 9323 15211
rect 8379 15147 8391 15199
rect 8443 15147 8515 15199
rect 8567 15147 8639 15199
rect 8691 15147 8763 15199
rect 8815 15147 8887 15199
rect 8939 15147 9011 15199
rect 9063 15147 9135 15199
rect 9187 15147 9259 15199
rect 9311 15147 9323 15199
rect 8379 15075 9323 15147
rect 8379 15023 8391 15075
rect 8443 15023 8515 15075
rect 8567 15023 8639 15075
rect 8691 15023 8763 15075
rect 8815 15023 8887 15075
rect 8939 15023 9011 15075
rect 9063 15023 9135 15075
rect 9187 15023 9259 15075
rect 9311 15023 9323 15075
rect 8379 14951 9323 15023
rect 8379 14899 8391 14951
rect 8443 14899 8515 14951
rect 8567 14899 8639 14951
rect 8691 14899 8763 14951
rect 8815 14899 8887 14951
rect 8939 14899 9011 14951
rect 9063 14899 9135 14951
rect 9187 14899 9259 14951
rect 9311 14899 9323 14951
rect 8379 14827 9323 14899
rect 8379 14775 8391 14827
rect 8443 14775 8515 14827
rect 8567 14775 8639 14827
rect 8691 14775 8763 14827
rect 8815 14775 8887 14827
rect 8939 14775 9011 14827
rect 9063 14775 9135 14827
rect 9187 14775 9259 14827
rect 9311 14775 9323 14827
rect 8379 14748 9323 14775
rect 8379 14703 8397 14748
rect 8453 14703 8539 14748
rect 8595 14703 8681 14748
rect 8737 14703 8823 14748
rect 8379 14651 8391 14703
rect 8453 14692 8515 14703
rect 8595 14692 8639 14703
rect 8737 14692 8763 14703
rect 8443 14651 8515 14692
rect 8567 14651 8639 14692
rect 8691 14651 8763 14692
rect 8815 14692 8823 14703
rect 8879 14703 8965 14748
rect 9021 14703 9107 14748
rect 9163 14703 9249 14748
rect 9305 14703 9323 14748
rect 8879 14692 8887 14703
rect 8815 14651 8887 14692
rect 8939 14692 8965 14703
rect 9063 14692 9107 14703
rect 9187 14692 9249 14703
rect 8939 14651 9011 14692
rect 9063 14651 9135 14692
rect 9187 14651 9259 14692
rect 9311 14651 9323 14703
rect 8379 14606 9323 14651
rect 8379 14579 8397 14606
rect 8453 14579 8539 14606
rect 8595 14579 8681 14606
rect 8737 14579 8823 14606
rect 8379 14527 8391 14579
rect 8453 14550 8515 14579
rect 8595 14550 8639 14579
rect 8737 14550 8763 14579
rect 8443 14527 8515 14550
rect 8567 14527 8639 14550
rect 8691 14527 8763 14550
rect 8815 14550 8823 14579
rect 8879 14579 8965 14606
rect 9021 14579 9107 14606
rect 9163 14579 9249 14606
rect 9305 14579 9323 14606
rect 8879 14550 8887 14579
rect 8815 14527 8887 14550
rect 8939 14550 8965 14579
rect 9063 14550 9107 14579
rect 9187 14550 9249 14579
rect 8939 14527 9011 14550
rect 9063 14527 9135 14550
rect 9187 14527 9259 14550
rect 9311 14527 9323 14579
rect 8379 14464 9323 14527
rect 8379 14455 8397 14464
rect 8453 14455 8539 14464
rect 8595 14455 8681 14464
rect 8737 14455 8823 14464
rect 8379 14403 8391 14455
rect 8453 14408 8515 14455
rect 8595 14408 8639 14455
rect 8737 14408 8763 14455
rect 8443 14403 8515 14408
rect 8567 14403 8639 14408
rect 8691 14403 8763 14408
rect 8815 14408 8823 14455
rect 8879 14455 8965 14464
rect 9021 14455 9107 14464
rect 9163 14455 9249 14464
rect 9305 14455 9323 14464
rect 8879 14408 8887 14455
rect 8815 14403 8887 14408
rect 8939 14408 8965 14455
rect 9063 14408 9107 14455
rect 9187 14408 9249 14455
rect 8939 14403 9011 14408
rect 9063 14403 9135 14408
rect 9187 14403 9259 14408
rect 9311 14403 9323 14455
rect 8379 14391 9323 14403
rect 10145 15199 11089 15211
rect 10145 15147 10157 15199
rect 10209 15147 10281 15199
rect 10333 15147 10405 15199
rect 10457 15147 10529 15199
rect 10581 15147 10653 15199
rect 10705 15147 10777 15199
rect 10829 15147 10901 15199
rect 10953 15147 11025 15199
rect 11077 15147 11089 15199
rect 10145 15075 11089 15147
rect 10145 15023 10157 15075
rect 10209 15023 10281 15075
rect 10333 15023 10405 15075
rect 10457 15023 10529 15075
rect 10581 15023 10653 15075
rect 10705 15023 10777 15075
rect 10829 15023 10901 15075
rect 10953 15023 11025 15075
rect 11077 15023 11089 15075
rect 10145 14951 11089 15023
rect 10145 14899 10157 14951
rect 10209 14899 10281 14951
rect 10333 14899 10405 14951
rect 10457 14899 10529 14951
rect 10581 14899 10653 14951
rect 10705 14899 10777 14951
rect 10829 14899 10901 14951
rect 10953 14899 11025 14951
rect 11077 14899 11089 14951
rect 10145 14827 11089 14899
rect 10145 14775 10157 14827
rect 10209 14775 10281 14827
rect 10333 14775 10405 14827
rect 10457 14775 10529 14827
rect 10581 14775 10653 14827
rect 10705 14775 10777 14827
rect 10829 14775 10901 14827
rect 10953 14775 11025 14827
rect 11077 14775 11089 14827
rect 10145 14748 11089 14775
rect 10145 14703 10163 14748
rect 10219 14703 10305 14748
rect 10361 14703 10447 14748
rect 10503 14703 10589 14748
rect 10145 14651 10157 14703
rect 10219 14692 10281 14703
rect 10361 14692 10405 14703
rect 10503 14692 10529 14703
rect 10209 14651 10281 14692
rect 10333 14651 10405 14692
rect 10457 14651 10529 14692
rect 10581 14692 10589 14703
rect 10645 14703 10731 14748
rect 10787 14703 10873 14748
rect 10929 14703 11015 14748
rect 11071 14703 11089 14748
rect 10645 14692 10653 14703
rect 10581 14651 10653 14692
rect 10705 14692 10731 14703
rect 10829 14692 10873 14703
rect 10953 14692 11015 14703
rect 10705 14651 10777 14692
rect 10829 14651 10901 14692
rect 10953 14651 11025 14692
rect 11077 14651 11089 14703
rect 10145 14606 11089 14651
rect 10145 14579 10163 14606
rect 10219 14579 10305 14606
rect 10361 14579 10447 14606
rect 10503 14579 10589 14606
rect 10145 14527 10157 14579
rect 10219 14550 10281 14579
rect 10361 14550 10405 14579
rect 10503 14550 10529 14579
rect 10209 14527 10281 14550
rect 10333 14527 10405 14550
rect 10457 14527 10529 14550
rect 10581 14550 10589 14579
rect 10645 14579 10731 14606
rect 10787 14579 10873 14606
rect 10929 14579 11015 14606
rect 11071 14579 11089 14606
rect 10645 14550 10653 14579
rect 10581 14527 10653 14550
rect 10705 14550 10731 14579
rect 10829 14550 10873 14579
rect 10953 14550 11015 14579
rect 10705 14527 10777 14550
rect 10829 14527 10901 14550
rect 10953 14527 11025 14550
rect 11077 14527 11089 14579
rect 10145 14464 11089 14527
rect 10145 14455 10163 14464
rect 10219 14455 10305 14464
rect 10361 14455 10447 14464
rect 10503 14455 10589 14464
rect 10145 14403 10157 14455
rect 10219 14408 10281 14455
rect 10361 14408 10405 14455
rect 10503 14408 10529 14455
rect 10209 14403 10281 14408
rect 10333 14403 10405 14408
rect 10457 14403 10529 14408
rect 10581 14408 10589 14455
rect 10645 14455 10731 14464
rect 10787 14455 10873 14464
rect 10929 14455 11015 14464
rect 11071 14455 11089 14464
rect 10645 14408 10653 14455
rect 10581 14403 10653 14408
rect 10705 14408 10731 14455
rect 10829 14408 10873 14455
rect 10953 14408 11015 14455
rect 10705 14403 10777 14408
rect 10829 14403 10901 14408
rect 10953 14403 11025 14408
rect 11077 14403 11089 14455
rect 10145 14391 11089 14403
rect 11545 15183 11945 15250
rect 11545 15131 11595 15183
rect 11647 15131 11719 15183
rect 11771 15131 11843 15183
rect 11895 15131 11945 15183
rect 11545 15059 11945 15131
rect 11545 15007 11595 15059
rect 11647 15007 11719 15059
rect 11771 15007 11843 15059
rect 11895 15007 11945 15059
rect 11545 14935 11945 15007
rect 11545 14883 11595 14935
rect 11647 14883 11719 14935
rect 11771 14883 11843 14935
rect 11895 14883 11945 14935
rect 11545 14811 11945 14883
rect 11545 14759 11595 14811
rect 11647 14759 11719 14811
rect 11771 14759 11843 14811
rect 11895 14759 11945 14811
rect 11545 14755 11945 14759
rect 11545 14699 11575 14755
rect 11631 14699 11717 14755
rect 11773 14699 11859 14755
rect 11915 14699 11945 14755
rect 11545 14687 11945 14699
rect 11545 14635 11595 14687
rect 11647 14635 11719 14687
rect 11771 14635 11843 14687
rect 11895 14635 11945 14687
rect 11545 14613 11945 14635
rect 11545 14557 11575 14613
rect 11631 14557 11717 14613
rect 11773 14557 11859 14613
rect 11915 14557 11945 14613
rect 11545 14471 11945 14557
rect 11545 14415 11575 14471
rect 11631 14415 11717 14471
rect 11773 14415 11859 14471
rect 11915 14415 11945 14471
rect 416 14273 446 14329
rect 502 14273 588 14329
rect 644 14273 730 14329
rect 786 14273 816 14329
rect 416 14187 816 14273
rect 416 14131 446 14187
rect 502 14131 588 14187
rect 644 14131 730 14187
rect 786 14131 816 14187
rect 416 14045 816 14131
rect 416 13989 446 14045
rect 502 13989 588 14045
rect 644 13989 730 14045
rect 786 13989 816 14045
rect 416 13903 816 13989
rect 416 13847 446 13903
rect 502 13847 588 13903
rect 644 13847 730 13903
rect 786 13847 816 13903
rect 416 13761 816 13847
rect 416 13705 446 13761
rect 502 13705 588 13761
rect 644 13705 730 13761
rect 786 13705 816 13761
rect 416 13619 816 13705
rect 416 13563 446 13619
rect 502 13563 588 13619
rect 644 13563 730 13619
rect 786 13563 816 13619
rect 416 13477 816 13563
rect 416 13421 446 13477
rect 502 13421 588 13477
rect 644 13421 730 13477
rect 786 13421 816 13477
rect 416 13388 816 13421
rect 11545 14329 11945 14415
rect 11545 14273 11575 14329
rect 11631 14273 11717 14329
rect 11773 14273 11859 14329
rect 11915 14273 11945 14329
rect 11545 14187 11945 14273
rect 11545 14131 11575 14187
rect 11631 14131 11717 14187
rect 11773 14131 11859 14187
rect 11915 14131 11945 14187
rect 11545 14045 11945 14131
rect 11545 13989 11575 14045
rect 11631 13989 11717 14045
rect 11773 13989 11859 14045
rect 11915 13989 11945 14045
rect 11545 13903 11945 13989
rect 11545 13847 11575 13903
rect 11631 13847 11717 13903
rect 11773 13847 11859 13903
rect 11915 13847 11945 13903
rect 11545 13761 11945 13847
rect 11545 13705 11575 13761
rect 11631 13705 11717 13761
rect 11773 13705 11859 13761
rect 11915 13705 11945 13761
rect 11545 13619 11945 13705
rect 11545 13563 11575 13619
rect 11631 13563 11717 13619
rect 11773 13563 11859 13619
rect 11915 13563 11945 13619
rect 11545 13477 11945 13563
rect 11545 13421 11575 13477
rect 11631 13421 11717 13477
rect 11773 13421 11859 13477
rect 11915 13421 11945 13477
rect 11545 13388 11945 13421
rect 428 13148 816 13188
rect 428 13092 452 13148
rect 508 13109 594 13148
rect 650 13109 736 13148
rect 524 13092 594 13109
rect 650 13092 720 13109
rect 792 13092 816 13148
rect 428 13057 472 13092
rect 524 13057 596 13092
rect 648 13057 720 13092
rect 772 13057 816 13092
rect 428 13006 816 13057
rect 428 12950 452 13006
rect 508 12985 594 13006
rect 650 12985 736 13006
rect 524 12950 594 12985
rect 650 12950 720 12985
rect 792 12950 816 13006
rect 428 12933 472 12950
rect 524 12933 596 12950
rect 648 12933 720 12950
rect 772 12933 816 12950
rect 428 12864 816 12933
rect 428 12808 452 12864
rect 508 12861 594 12864
rect 650 12861 736 12864
rect 524 12809 594 12861
rect 650 12809 720 12861
rect 508 12808 594 12809
rect 650 12808 736 12809
rect 792 12808 816 12864
rect 428 12737 816 12808
rect 428 12722 472 12737
rect 524 12722 596 12737
rect 648 12722 720 12737
rect 772 12722 816 12737
rect 428 12666 452 12722
rect 524 12685 594 12722
rect 650 12685 720 12722
rect 508 12666 594 12685
rect 650 12666 736 12685
rect 792 12666 816 12722
rect 428 12613 816 12666
rect 428 12580 472 12613
rect 524 12580 596 12613
rect 648 12580 720 12613
rect 772 12580 816 12613
rect 428 12524 452 12580
rect 524 12561 594 12580
rect 650 12561 720 12580
rect 508 12524 594 12561
rect 650 12524 736 12561
rect 792 12524 816 12580
rect 428 12489 816 12524
rect 428 12438 472 12489
rect 524 12438 596 12489
rect 648 12438 720 12489
rect 772 12438 816 12489
rect 428 12382 452 12438
rect 524 12437 594 12438
rect 650 12437 720 12438
rect 508 12382 594 12437
rect 650 12382 736 12437
rect 792 12382 816 12438
rect 428 12365 816 12382
rect 428 12313 472 12365
rect 524 12313 596 12365
rect 648 12313 720 12365
rect 772 12313 816 12365
rect 428 12296 816 12313
rect 428 12240 452 12296
rect 508 12241 594 12296
rect 650 12241 736 12296
rect 524 12240 594 12241
rect 650 12240 720 12241
rect 792 12240 816 12296
rect 428 12189 472 12240
rect 524 12189 596 12240
rect 648 12189 720 12240
rect 772 12189 816 12240
rect 428 12154 816 12189
rect 428 12098 452 12154
rect 508 12117 594 12154
rect 650 12117 736 12154
rect 524 12098 594 12117
rect 650 12098 720 12117
rect 792 12098 816 12154
rect 428 12065 472 12098
rect 524 12065 596 12098
rect 648 12065 720 12098
rect 772 12065 816 12098
rect 428 12012 816 12065
rect 428 11956 452 12012
rect 508 11993 594 12012
rect 650 11993 736 12012
rect 524 11956 594 11993
rect 650 11956 720 11993
rect 792 11956 816 12012
rect 428 11941 472 11956
rect 524 11941 596 11956
rect 648 11941 720 11956
rect 772 11941 816 11956
rect 428 11870 816 11941
rect 428 11814 452 11870
rect 508 11869 594 11870
rect 650 11869 736 11870
rect 524 11817 594 11869
rect 650 11817 720 11869
rect 508 11814 594 11817
rect 650 11814 736 11817
rect 792 11814 816 11870
rect 428 11745 816 11814
rect 428 11728 472 11745
rect 524 11728 596 11745
rect 648 11728 720 11745
rect 772 11728 816 11745
rect 428 11672 452 11728
rect 524 11693 594 11728
rect 650 11693 720 11728
rect 508 11672 594 11693
rect 650 11672 736 11693
rect 792 11672 816 11728
rect 428 11621 816 11672
rect 428 11586 472 11621
rect 524 11586 596 11621
rect 648 11586 720 11621
rect 772 11586 816 11621
rect 428 11530 452 11586
rect 524 11569 594 11586
rect 650 11569 720 11586
rect 508 11530 594 11569
rect 650 11530 736 11569
rect 792 11530 816 11586
rect 428 11472 816 11530
rect 11557 13148 11945 13188
rect 11557 13092 11581 13148
rect 11637 13109 11723 13148
rect 11779 13109 11865 13148
rect 11653 13092 11723 13109
rect 11779 13092 11849 13109
rect 11921 13092 11945 13148
rect 11557 13057 11601 13092
rect 11653 13057 11725 13092
rect 11777 13057 11849 13092
rect 11901 13057 11945 13092
rect 11557 13006 11945 13057
rect 11557 12950 11581 13006
rect 11637 12985 11723 13006
rect 11779 12985 11865 13006
rect 11653 12950 11723 12985
rect 11779 12950 11849 12985
rect 11921 12950 11945 13006
rect 11557 12933 11601 12950
rect 11653 12933 11725 12950
rect 11777 12933 11849 12950
rect 11901 12933 11945 12950
rect 11557 12864 11945 12933
rect 11557 12808 11581 12864
rect 11637 12861 11723 12864
rect 11779 12861 11865 12864
rect 11653 12809 11723 12861
rect 11779 12809 11849 12861
rect 11637 12808 11723 12809
rect 11779 12808 11865 12809
rect 11921 12808 11945 12864
rect 11557 12737 11945 12808
rect 11557 12722 11601 12737
rect 11653 12722 11725 12737
rect 11777 12722 11849 12737
rect 11901 12722 11945 12737
rect 11557 12666 11581 12722
rect 11653 12685 11723 12722
rect 11779 12685 11849 12722
rect 11637 12666 11723 12685
rect 11779 12666 11865 12685
rect 11921 12666 11945 12722
rect 11557 12613 11945 12666
rect 11557 12580 11601 12613
rect 11653 12580 11725 12613
rect 11777 12580 11849 12613
rect 11901 12580 11945 12613
rect 11557 12524 11581 12580
rect 11653 12561 11723 12580
rect 11779 12561 11849 12580
rect 11637 12524 11723 12561
rect 11779 12524 11865 12561
rect 11921 12524 11945 12580
rect 11557 12489 11945 12524
rect 11557 12438 11601 12489
rect 11653 12438 11725 12489
rect 11777 12438 11849 12489
rect 11901 12438 11945 12489
rect 11557 12382 11581 12438
rect 11653 12437 11723 12438
rect 11779 12437 11849 12438
rect 11637 12382 11723 12437
rect 11779 12382 11865 12437
rect 11921 12382 11945 12438
rect 11557 12365 11945 12382
rect 11557 12313 11601 12365
rect 11653 12313 11725 12365
rect 11777 12313 11849 12365
rect 11901 12313 11945 12365
rect 11557 12296 11945 12313
rect 11557 12240 11581 12296
rect 11637 12241 11723 12296
rect 11779 12241 11865 12296
rect 11653 12240 11723 12241
rect 11779 12240 11849 12241
rect 11921 12240 11945 12296
rect 11557 12189 11601 12240
rect 11653 12189 11725 12240
rect 11777 12189 11849 12240
rect 11901 12189 11945 12240
rect 11557 12154 11945 12189
rect 11557 12098 11581 12154
rect 11637 12117 11723 12154
rect 11779 12117 11865 12154
rect 11653 12098 11723 12117
rect 11779 12098 11849 12117
rect 11921 12098 11945 12154
rect 11557 12065 11601 12098
rect 11653 12065 11725 12098
rect 11777 12065 11849 12098
rect 11901 12065 11945 12098
rect 11557 12012 11945 12065
rect 11557 11956 11581 12012
rect 11637 11993 11723 12012
rect 11779 11993 11865 12012
rect 11653 11956 11723 11993
rect 11779 11956 11849 11993
rect 11921 11956 11945 12012
rect 11557 11941 11601 11956
rect 11653 11941 11725 11956
rect 11777 11941 11849 11956
rect 11901 11941 11945 11956
rect 11557 11870 11945 11941
rect 11557 11814 11581 11870
rect 11637 11869 11723 11870
rect 11779 11869 11865 11870
rect 11653 11817 11723 11869
rect 11779 11817 11849 11869
rect 11637 11814 11723 11817
rect 11779 11814 11865 11817
rect 11921 11814 11945 11870
rect 11557 11745 11945 11814
rect 11557 11728 11601 11745
rect 11653 11728 11725 11745
rect 11777 11728 11849 11745
rect 11901 11728 11945 11745
rect 11557 11672 11581 11728
rect 11653 11693 11723 11728
rect 11779 11693 11849 11728
rect 11637 11672 11723 11693
rect 11779 11672 11865 11693
rect 11921 11672 11945 11728
rect 11557 11621 11945 11672
rect 11557 11586 11601 11621
rect 11653 11586 11725 11621
rect 11777 11586 11849 11621
rect 11901 11586 11945 11621
rect 11557 11530 11581 11586
rect 11653 11569 11723 11586
rect 11779 11569 11849 11586
rect 11637 11530 11723 11569
rect 11779 11530 11865 11569
rect 11921 11530 11945 11586
rect 11557 11472 11945 11530
rect 428 10887 1009 10972
rect 428 10861 471 10887
rect 527 10861 613 10887
rect 669 10861 1009 10887
rect 428 10289 440 10861
rect 700 10289 1009 10861
rect 428 10263 471 10289
rect 527 10263 613 10289
rect 669 10263 1009 10289
rect 428 10188 1009 10263
rect 11373 10887 11954 10972
rect 11373 10861 11713 10887
rect 11769 10861 11855 10887
rect 11911 10861 11954 10887
rect 11373 10289 11682 10861
rect 11942 10289 11954 10861
rect 11373 10263 11713 10289
rect 11769 10263 11855 10289
rect 11911 10263 11954 10289
rect 11373 10188 11954 10263
rect 428 9922 1009 9988
rect 428 9866 471 9922
rect 527 9866 613 9922
rect 669 9866 1009 9922
rect 428 9852 1009 9866
rect 428 7096 440 9852
rect 700 7096 1009 9852
rect 428 7082 1009 7096
rect 428 7026 471 7082
rect 527 7026 613 7082
rect 669 7026 1009 7082
rect 428 6988 1009 7026
rect 11373 9922 11954 9988
rect 11373 9866 11713 9922
rect 11769 9866 11855 9922
rect 11911 9866 11954 9922
rect 11373 9852 11954 9866
rect 11373 7096 11682 9852
rect 11942 7096 11954 9852
rect 11373 7082 11954 7096
rect 11373 7026 11713 7082
rect 11769 7026 11855 7082
rect 11911 7026 11954 7082
rect 11373 6988 11954 7026
rect 428 6740 1009 6788
rect 428 6684 471 6740
rect 527 6684 613 6740
rect 669 6684 1009 6740
rect 428 6682 1009 6684
rect 428 3926 440 6682
rect 700 3926 1009 6682
rect 428 3900 1009 3926
rect 428 3844 471 3900
rect 527 3844 613 3900
rect 669 3844 1009 3900
rect 428 3788 1009 3844
rect 11373 6740 11954 6788
rect 11373 6684 11713 6740
rect 11769 6684 11855 6740
rect 11911 6684 11954 6740
rect 11373 6682 11954 6684
rect 11373 3926 11682 6682
rect 11942 3926 11954 6682
rect 11373 3900 11954 3926
rect 11373 3844 11713 3900
rect 11769 3844 11855 3900
rect 11911 3844 11954 3900
rect 11373 3788 11954 3844
rect 428 3522 1009 3588
rect 428 3505 471 3522
rect 527 3505 613 3522
rect 669 3505 1009 3522
rect 428 3037 440 3505
rect 700 3037 1009 3505
rect 428 2972 1009 3037
rect 11373 3522 11954 3588
rect 11373 3505 11713 3522
rect 11769 3505 11855 3522
rect 11911 3505 11954 3522
rect 11373 3037 11682 3505
rect 11942 3037 11954 3505
rect 11373 2972 11954 3037
rect 428 2402 816 2414
rect 428 2350 472 2402
rect 524 2350 596 2402
rect 648 2350 720 2402
rect 772 2350 816 2402
rect 428 2317 816 2350
rect 428 2261 452 2317
rect 508 2278 594 2317
rect 650 2278 736 2317
rect 524 2261 594 2278
rect 650 2261 720 2278
rect 792 2261 816 2317
rect 428 2226 472 2261
rect 524 2226 596 2261
rect 648 2226 720 2261
rect 772 2226 816 2261
rect 428 2175 816 2226
rect 428 2119 452 2175
rect 508 2154 594 2175
rect 650 2154 736 2175
rect 524 2119 594 2154
rect 650 2119 720 2154
rect 792 2119 816 2175
rect 428 2102 472 2119
rect 524 2102 596 2119
rect 648 2102 720 2119
rect 772 2102 816 2119
rect 428 2033 816 2102
rect 428 1977 452 2033
rect 508 2030 594 2033
rect 650 2030 736 2033
rect 524 1978 594 2030
rect 650 1978 720 2030
rect 508 1977 594 1978
rect 650 1977 736 1978
rect 792 1977 816 2033
rect 428 1906 816 1977
rect 428 1891 472 1906
rect 524 1891 596 1906
rect 648 1891 720 1906
rect 772 1891 816 1906
rect 428 1835 452 1891
rect 524 1854 594 1891
rect 650 1854 720 1891
rect 508 1835 594 1854
rect 650 1835 736 1854
rect 792 1835 816 1891
rect 428 1782 816 1835
rect 428 1749 472 1782
rect 524 1749 596 1782
rect 648 1749 720 1782
rect 772 1749 816 1782
rect 428 1693 452 1749
rect 524 1730 594 1749
rect 650 1730 720 1749
rect 508 1693 594 1730
rect 650 1693 736 1730
rect 792 1693 816 1749
rect 428 1658 816 1693
rect 428 1607 472 1658
rect 524 1607 596 1658
rect 648 1607 720 1658
rect 772 1607 816 1658
rect 428 1551 452 1607
rect 524 1606 594 1607
rect 650 1606 720 1607
rect 508 1551 594 1606
rect 650 1551 736 1606
rect 792 1551 816 1607
rect 428 1534 816 1551
rect 428 1482 472 1534
rect 524 1482 596 1534
rect 648 1482 720 1534
rect 772 1482 816 1534
rect 428 1465 816 1482
rect 428 1409 452 1465
rect 508 1410 594 1465
rect 650 1410 736 1465
rect 524 1409 594 1410
rect 650 1409 720 1410
rect 792 1409 816 1465
rect 428 1358 472 1409
rect 524 1358 596 1409
rect 648 1358 720 1409
rect 772 1358 816 1409
rect 428 1323 816 1358
rect 428 1267 452 1323
rect 508 1286 594 1323
rect 650 1286 736 1323
rect 524 1267 594 1286
rect 650 1267 720 1286
rect 792 1267 816 1323
rect 428 1234 472 1267
rect 524 1234 596 1267
rect 648 1234 720 1267
rect 772 1234 816 1267
rect 428 1181 816 1234
rect 428 1125 452 1181
rect 508 1162 594 1181
rect 650 1162 736 1181
rect 524 1125 594 1162
rect 650 1125 720 1162
rect 792 1125 816 1181
rect 428 1110 472 1125
rect 524 1110 596 1125
rect 648 1110 720 1125
rect 772 1110 816 1125
rect 428 1039 816 1110
rect 428 983 452 1039
rect 508 1038 594 1039
rect 650 1038 736 1039
rect 524 986 594 1038
rect 650 986 720 1038
rect 508 983 594 986
rect 650 983 736 986
rect 792 983 816 1039
rect 428 914 816 983
rect 428 897 472 914
rect 524 897 596 914
rect 648 897 720 914
rect 772 897 816 914
rect 428 841 452 897
rect 524 862 594 897
rect 650 862 720 897
rect 508 841 594 862
rect 650 841 736 862
rect 792 841 816 897
rect 428 790 816 841
rect 428 755 472 790
rect 524 755 596 790
rect 648 755 720 790
rect 772 755 816 790
rect 428 699 452 755
rect 524 738 594 755
rect 650 738 720 755
rect 508 699 594 738
rect 650 699 736 738
rect 792 699 816 755
rect 428 666 816 699
rect 428 614 472 666
rect 524 614 596 666
rect 648 614 720 666
rect 772 614 816 666
rect 428 602 816 614
rect 11557 2402 11945 2414
rect 11557 2350 11601 2402
rect 11653 2350 11725 2402
rect 11777 2350 11849 2402
rect 11901 2350 11945 2402
rect 11557 2317 11945 2350
rect 11557 2261 11581 2317
rect 11637 2278 11723 2317
rect 11779 2278 11865 2317
rect 11653 2261 11723 2278
rect 11779 2261 11849 2278
rect 11921 2261 11945 2317
rect 11557 2226 11601 2261
rect 11653 2226 11725 2261
rect 11777 2226 11849 2261
rect 11901 2226 11945 2261
rect 11557 2175 11945 2226
rect 11557 2119 11581 2175
rect 11637 2154 11723 2175
rect 11779 2154 11865 2175
rect 11653 2119 11723 2154
rect 11779 2119 11849 2154
rect 11921 2119 11945 2175
rect 11557 2102 11601 2119
rect 11653 2102 11725 2119
rect 11777 2102 11849 2119
rect 11901 2102 11945 2119
rect 11557 2033 11945 2102
rect 11557 1977 11581 2033
rect 11637 2030 11723 2033
rect 11779 2030 11865 2033
rect 11653 1978 11723 2030
rect 11779 1978 11849 2030
rect 11637 1977 11723 1978
rect 11779 1977 11865 1978
rect 11921 1977 11945 2033
rect 11557 1906 11945 1977
rect 11557 1891 11601 1906
rect 11653 1891 11725 1906
rect 11777 1891 11849 1906
rect 11901 1891 11945 1906
rect 11557 1835 11581 1891
rect 11653 1854 11723 1891
rect 11779 1854 11849 1891
rect 11637 1835 11723 1854
rect 11779 1835 11865 1854
rect 11921 1835 11945 1891
rect 11557 1782 11945 1835
rect 11557 1749 11601 1782
rect 11653 1749 11725 1782
rect 11777 1749 11849 1782
rect 11901 1749 11945 1782
rect 11557 1693 11581 1749
rect 11653 1730 11723 1749
rect 11779 1730 11849 1749
rect 11637 1693 11723 1730
rect 11779 1693 11865 1730
rect 11921 1693 11945 1749
rect 11557 1658 11945 1693
rect 11557 1607 11601 1658
rect 11653 1607 11725 1658
rect 11777 1607 11849 1658
rect 11901 1607 11945 1658
rect 11557 1551 11581 1607
rect 11653 1606 11723 1607
rect 11779 1606 11849 1607
rect 11637 1551 11723 1606
rect 11779 1551 11865 1606
rect 11921 1551 11945 1607
rect 11557 1534 11945 1551
rect 11557 1482 11601 1534
rect 11653 1482 11725 1534
rect 11777 1482 11849 1534
rect 11901 1482 11945 1534
rect 11557 1465 11945 1482
rect 11557 1409 11581 1465
rect 11637 1410 11723 1465
rect 11779 1410 11865 1465
rect 11653 1409 11723 1410
rect 11779 1409 11849 1410
rect 11921 1409 11945 1465
rect 11557 1358 11601 1409
rect 11653 1358 11725 1409
rect 11777 1358 11849 1409
rect 11901 1358 11945 1409
rect 11557 1323 11945 1358
rect 11557 1267 11581 1323
rect 11637 1286 11723 1323
rect 11779 1286 11865 1323
rect 11653 1267 11723 1286
rect 11779 1267 11849 1286
rect 11921 1267 11945 1323
rect 11557 1234 11601 1267
rect 11653 1234 11725 1267
rect 11777 1234 11849 1267
rect 11901 1234 11945 1267
rect 11557 1181 11945 1234
rect 11557 1125 11581 1181
rect 11637 1162 11723 1181
rect 11779 1162 11865 1181
rect 11653 1125 11723 1162
rect 11779 1125 11849 1162
rect 11921 1125 11945 1181
rect 11557 1110 11601 1125
rect 11653 1110 11725 1125
rect 11777 1110 11849 1125
rect 11901 1110 11945 1125
rect 11557 1039 11945 1110
rect 11557 983 11581 1039
rect 11637 1038 11723 1039
rect 11779 1038 11865 1039
rect 11653 986 11723 1038
rect 11779 986 11849 1038
rect 11637 983 11723 986
rect 11779 983 11865 986
rect 11921 983 11945 1039
rect 11557 914 11945 983
rect 11557 897 11601 914
rect 11653 897 11725 914
rect 11777 897 11849 914
rect 11901 897 11945 914
rect 11557 841 11581 897
rect 11653 862 11723 897
rect 11779 862 11849 897
rect 11637 841 11723 862
rect 11779 841 11865 862
rect 11921 841 11945 897
rect 11557 790 11945 841
rect 11557 755 11601 790
rect 11653 755 11725 790
rect 11777 755 11849 790
rect 11901 755 11945 790
rect 11557 699 11581 755
rect 11653 738 11723 755
rect 11779 738 11849 755
rect 11637 699 11723 738
rect 11779 699 11865 738
rect 11921 699 11945 755
rect 11557 666 11945 699
rect 11557 614 11601 666
rect 11653 614 11725 666
rect 11777 614 11849 666
rect 11901 614 11945 666
rect 11557 602 11945 614
rect 12860 356 13078 366
rect -708 298 -528 302
rect 12860 300 12870 356
rect 12926 339 13012 356
rect 13068 300 13078 356
rect -727 290 -509 298
rect -727 288 -696 290
rect -540 288 -509 290
rect -727 232 -717 288
rect -519 232 -509 288
rect -727 146 -696 232
rect -540 146 -509 232
rect -727 90 -717 146
rect -519 90 -509 146
rect -727 4 -696 90
rect -540 4 -509 90
rect -727 -52 -717 4
rect -519 -52 -509 4
rect -727 -138 -696 -52
rect -540 -138 -509 -52
rect -727 -194 -717 -138
rect -519 -194 -509 -138
rect -727 -280 -696 -194
rect -540 -280 -509 -194
rect -727 -336 -717 -280
rect -519 -336 -509 -280
rect -727 -422 -696 -336
rect -540 -422 -509 -336
rect -727 -478 -717 -422
rect -519 -478 -509 -422
rect -727 -564 -696 -478
rect -540 -564 -509 -478
rect -727 -620 -717 -564
rect -519 -620 -509 -564
rect -727 -706 -696 -620
rect -540 -706 -509 -620
rect -727 -762 -717 -706
rect -519 -762 -509 -706
rect -727 -848 -696 -762
rect -540 -848 -509 -762
rect -727 -904 -717 -848
rect -519 -904 -509 -848
rect -727 -906 -696 -904
rect -540 -906 -509 -904
rect -727 -914 -509 -906
rect 12860 214 12891 300
rect 13047 214 13078 300
rect 12860 158 12870 214
rect 13068 158 13078 214
rect 12860 72 12891 158
rect 13047 72 13078 158
rect 12860 16 12870 72
rect 13068 16 13078 72
rect 12860 -70 12891 16
rect 13047 -70 13078 16
rect 12860 -126 12870 -70
rect 13068 -126 13078 -70
rect 12860 -212 12891 -126
rect 13047 -212 13078 -126
rect 12860 -268 12870 -212
rect 13068 -268 13078 -212
rect 12860 -354 12891 -268
rect 13047 -354 13078 -268
rect 12860 -410 12870 -354
rect 13068 -410 13078 -354
rect 12860 -496 12891 -410
rect 13047 -496 13078 -410
rect 12860 -552 12870 -496
rect 13068 -552 13078 -496
rect 12860 -638 12891 -552
rect 13047 -638 13078 -552
rect 12860 -694 12870 -638
rect 13068 -694 13078 -638
rect 12860 -780 12891 -694
rect 13047 -780 13078 -694
rect 12860 -836 12870 -780
rect 13068 -836 13078 -780
rect -708 -918 -528 -914
rect 12860 -922 12891 -836
rect 13047 -922 13078 -836
rect 12860 -978 12870 -922
rect 12926 -978 13012 -961
rect 13068 -978 13078 -922
rect 12860 -988 13078 -978
<< via2 >>
rect -684 14708 -628 14755
rect -542 14708 -486 14755
rect -684 14699 -667 14708
rect -667 14699 -628 14708
rect -542 14699 -503 14708
rect -503 14699 -486 14708
rect -684 14600 -628 14613
rect -542 14600 -486 14613
rect -684 14557 -667 14600
rect -667 14557 -628 14600
rect -542 14557 -503 14600
rect -503 14557 -486 14600
rect -684 14440 -667 14471
rect -667 14440 -628 14471
rect -542 14440 -503 14471
rect -503 14440 -486 14471
rect -684 14415 -628 14440
rect -542 14415 -486 14440
rect -684 14276 -628 14329
rect -542 14276 -486 14329
rect -684 14273 -667 14276
rect -667 14273 -628 14276
rect -542 14273 -503 14276
rect -503 14273 -486 14276
rect -684 14168 -628 14187
rect -542 14168 -486 14187
rect -684 14131 -667 14168
rect -667 14131 -628 14168
rect -542 14131 -503 14168
rect -503 14131 -486 14168
rect -684 14008 -667 14045
rect -667 14008 -628 14045
rect -542 14008 -503 14045
rect -503 14008 -486 14045
rect -684 13989 -628 14008
rect -542 13989 -486 14008
rect -684 13900 -667 13903
rect -667 13900 -628 13903
rect -542 13900 -503 13903
rect -503 13900 -486 13903
rect -684 13847 -628 13900
rect -542 13847 -486 13900
rect -684 13736 -628 13761
rect -542 13736 -486 13761
rect -684 13705 -667 13736
rect -667 13705 -628 13736
rect -542 13705 -503 13736
rect -503 13705 -486 13736
rect -684 13576 -667 13619
rect -667 13576 -628 13619
rect -542 13576 -503 13619
rect -503 13576 -486 13619
rect -684 13563 -628 13576
rect -542 13563 -486 13576
rect -684 13468 -667 13477
rect -667 13468 -628 13477
rect -542 13468 -503 13477
rect -503 13468 -486 13477
rect -684 13421 -628 13468
rect -542 13421 -486 13468
rect 446 14699 502 14755
rect 588 14699 644 14755
rect 730 14699 786 14755
rect 446 14557 502 14613
rect 588 14557 644 14613
rect 730 14557 786 14613
rect 446 14415 502 14471
rect 588 14415 644 14471
rect 730 14415 786 14471
rect 1322 14703 1378 14748
rect 1464 14703 1520 14748
rect 1606 14703 1662 14748
rect 1322 14692 1368 14703
rect 1368 14692 1378 14703
rect 1464 14692 1492 14703
rect 1492 14692 1520 14703
rect 1606 14692 1616 14703
rect 1616 14692 1662 14703
rect 1748 14692 1804 14748
rect 1890 14703 1946 14748
rect 2032 14703 2088 14748
rect 2174 14703 2230 14748
rect 1890 14692 1936 14703
rect 1936 14692 1946 14703
rect 2032 14692 2060 14703
rect 2060 14692 2088 14703
rect 2174 14692 2184 14703
rect 2184 14692 2230 14703
rect 1322 14579 1378 14606
rect 1464 14579 1520 14606
rect 1606 14579 1662 14606
rect 1322 14550 1368 14579
rect 1368 14550 1378 14579
rect 1464 14550 1492 14579
rect 1492 14550 1520 14579
rect 1606 14550 1616 14579
rect 1616 14550 1662 14579
rect 1748 14550 1804 14606
rect 1890 14579 1946 14606
rect 2032 14579 2088 14606
rect 2174 14579 2230 14606
rect 1890 14550 1936 14579
rect 1936 14550 1946 14579
rect 2032 14550 2060 14579
rect 2060 14550 2088 14579
rect 2174 14550 2184 14579
rect 2184 14550 2230 14579
rect 1322 14455 1378 14464
rect 1464 14455 1520 14464
rect 1606 14455 1662 14464
rect 1322 14408 1368 14455
rect 1368 14408 1378 14455
rect 1464 14408 1492 14455
rect 1492 14408 1520 14455
rect 1606 14408 1616 14455
rect 1616 14408 1662 14455
rect 1748 14408 1804 14464
rect 1890 14455 1946 14464
rect 2032 14455 2088 14464
rect 2174 14455 2230 14464
rect 1890 14408 1936 14455
rect 1936 14408 1946 14455
rect 2032 14408 2060 14455
rect 2060 14408 2088 14455
rect 2174 14408 2184 14455
rect 2184 14408 2230 14455
rect 3094 14703 3150 14748
rect 3236 14703 3292 14748
rect 3378 14703 3434 14748
rect 3094 14692 3140 14703
rect 3140 14692 3150 14703
rect 3236 14692 3264 14703
rect 3264 14692 3292 14703
rect 3378 14692 3388 14703
rect 3388 14692 3434 14703
rect 3520 14692 3576 14748
rect 3662 14703 3718 14748
rect 3804 14703 3860 14748
rect 3946 14703 4002 14748
rect 3662 14692 3708 14703
rect 3708 14692 3718 14703
rect 3804 14692 3832 14703
rect 3832 14692 3860 14703
rect 3946 14692 3956 14703
rect 3956 14692 4002 14703
rect 3094 14579 3150 14606
rect 3236 14579 3292 14606
rect 3378 14579 3434 14606
rect 3094 14550 3140 14579
rect 3140 14550 3150 14579
rect 3236 14550 3264 14579
rect 3264 14550 3292 14579
rect 3378 14550 3388 14579
rect 3388 14550 3434 14579
rect 3520 14550 3576 14606
rect 3662 14579 3718 14606
rect 3804 14579 3860 14606
rect 3946 14579 4002 14606
rect 3662 14550 3708 14579
rect 3708 14550 3718 14579
rect 3804 14550 3832 14579
rect 3832 14550 3860 14579
rect 3946 14550 3956 14579
rect 3956 14550 4002 14579
rect 3094 14455 3150 14464
rect 3236 14455 3292 14464
rect 3378 14455 3434 14464
rect 3094 14408 3140 14455
rect 3140 14408 3150 14455
rect 3236 14408 3264 14455
rect 3264 14408 3292 14455
rect 3378 14408 3388 14455
rect 3388 14408 3434 14455
rect 3520 14408 3576 14464
rect 3662 14455 3718 14464
rect 3804 14455 3860 14464
rect 3946 14455 4002 14464
rect 3662 14408 3708 14455
rect 3708 14408 3718 14455
rect 3804 14408 3832 14455
rect 3832 14408 3860 14455
rect 3946 14408 3956 14455
rect 3956 14408 4002 14455
rect 4859 14703 4915 14748
rect 5001 14703 5057 14748
rect 5143 14703 5199 14748
rect 4859 14692 4905 14703
rect 4905 14692 4915 14703
rect 5001 14692 5029 14703
rect 5029 14692 5057 14703
rect 5143 14692 5153 14703
rect 5153 14692 5199 14703
rect 5285 14692 5341 14748
rect 5427 14703 5483 14748
rect 5569 14703 5625 14748
rect 5711 14703 5767 14748
rect 5427 14692 5473 14703
rect 5473 14692 5483 14703
rect 5569 14692 5597 14703
rect 5597 14692 5625 14703
rect 5711 14692 5721 14703
rect 5721 14692 5767 14703
rect 4859 14579 4915 14606
rect 5001 14579 5057 14606
rect 5143 14579 5199 14606
rect 4859 14550 4905 14579
rect 4905 14550 4915 14579
rect 5001 14550 5029 14579
rect 5029 14550 5057 14579
rect 5143 14550 5153 14579
rect 5153 14550 5199 14579
rect 5285 14550 5341 14606
rect 5427 14579 5483 14606
rect 5569 14579 5625 14606
rect 5711 14579 5767 14606
rect 5427 14550 5473 14579
rect 5473 14550 5483 14579
rect 5569 14550 5597 14579
rect 5597 14550 5625 14579
rect 5711 14550 5721 14579
rect 5721 14550 5767 14579
rect 4859 14455 4915 14464
rect 5001 14455 5057 14464
rect 5143 14455 5199 14464
rect 4859 14408 4905 14455
rect 4905 14408 4915 14455
rect 5001 14408 5029 14455
rect 5029 14408 5057 14455
rect 5143 14408 5153 14455
rect 5153 14408 5199 14455
rect 5285 14408 5341 14464
rect 5427 14455 5483 14464
rect 5569 14455 5625 14464
rect 5711 14455 5767 14464
rect 5427 14408 5473 14455
rect 5473 14408 5483 14455
rect 5569 14408 5597 14455
rect 5597 14408 5625 14455
rect 5711 14408 5721 14455
rect 5721 14408 5767 14455
rect 6628 14703 6684 14748
rect 6770 14703 6826 14748
rect 6912 14703 6968 14748
rect 6628 14692 6674 14703
rect 6674 14692 6684 14703
rect 6770 14692 6798 14703
rect 6798 14692 6826 14703
rect 6912 14692 6922 14703
rect 6922 14692 6968 14703
rect 7054 14692 7110 14748
rect 7196 14703 7252 14748
rect 7338 14703 7394 14748
rect 7480 14703 7536 14748
rect 7196 14692 7242 14703
rect 7242 14692 7252 14703
rect 7338 14692 7366 14703
rect 7366 14692 7394 14703
rect 7480 14692 7490 14703
rect 7490 14692 7536 14703
rect 6628 14579 6684 14606
rect 6770 14579 6826 14606
rect 6912 14579 6968 14606
rect 6628 14550 6674 14579
rect 6674 14550 6684 14579
rect 6770 14550 6798 14579
rect 6798 14550 6826 14579
rect 6912 14550 6922 14579
rect 6922 14550 6968 14579
rect 7054 14550 7110 14606
rect 7196 14579 7252 14606
rect 7338 14579 7394 14606
rect 7480 14579 7536 14606
rect 7196 14550 7242 14579
rect 7242 14550 7252 14579
rect 7338 14550 7366 14579
rect 7366 14550 7394 14579
rect 7480 14550 7490 14579
rect 7490 14550 7536 14579
rect 6628 14455 6684 14464
rect 6770 14455 6826 14464
rect 6912 14455 6968 14464
rect 6628 14408 6674 14455
rect 6674 14408 6684 14455
rect 6770 14408 6798 14455
rect 6798 14408 6826 14455
rect 6912 14408 6922 14455
rect 6922 14408 6968 14455
rect 7054 14408 7110 14464
rect 7196 14455 7252 14464
rect 7338 14455 7394 14464
rect 7480 14455 7536 14464
rect 7196 14408 7242 14455
rect 7242 14408 7252 14455
rect 7338 14408 7366 14455
rect 7366 14408 7394 14455
rect 7480 14408 7490 14455
rect 7490 14408 7536 14455
rect 8397 14703 8453 14748
rect 8539 14703 8595 14748
rect 8681 14703 8737 14748
rect 8397 14692 8443 14703
rect 8443 14692 8453 14703
rect 8539 14692 8567 14703
rect 8567 14692 8595 14703
rect 8681 14692 8691 14703
rect 8691 14692 8737 14703
rect 8823 14692 8879 14748
rect 8965 14703 9021 14748
rect 9107 14703 9163 14748
rect 9249 14703 9305 14748
rect 8965 14692 9011 14703
rect 9011 14692 9021 14703
rect 9107 14692 9135 14703
rect 9135 14692 9163 14703
rect 9249 14692 9259 14703
rect 9259 14692 9305 14703
rect 8397 14579 8453 14606
rect 8539 14579 8595 14606
rect 8681 14579 8737 14606
rect 8397 14550 8443 14579
rect 8443 14550 8453 14579
rect 8539 14550 8567 14579
rect 8567 14550 8595 14579
rect 8681 14550 8691 14579
rect 8691 14550 8737 14579
rect 8823 14550 8879 14606
rect 8965 14579 9021 14606
rect 9107 14579 9163 14606
rect 9249 14579 9305 14606
rect 8965 14550 9011 14579
rect 9011 14550 9021 14579
rect 9107 14550 9135 14579
rect 9135 14550 9163 14579
rect 9249 14550 9259 14579
rect 9259 14550 9305 14579
rect 8397 14455 8453 14464
rect 8539 14455 8595 14464
rect 8681 14455 8737 14464
rect 8397 14408 8443 14455
rect 8443 14408 8453 14455
rect 8539 14408 8567 14455
rect 8567 14408 8595 14455
rect 8681 14408 8691 14455
rect 8691 14408 8737 14455
rect 8823 14408 8879 14464
rect 8965 14455 9021 14464
rect 9107 14455 9163 14464
rect 9249 14455 9305 14464
rect 8965 14408 9011 14455
rect 9011 14408 9021 14455
rect 9107 14408 9135 14455
rect 9135 14408 9163 14455
rect 9249 14408 9259 14455
rect 9259 14408 9305 14455
rect 10163 14703 10219 14748
rect 10305 14703 10361 14748
rect 10447 14703 10503 14748
rect 10163 14692 10209 14703
rect 10209 14692 10219 14703
rect 10305 14692 10333 14703
rect 10333 14692 10361 14703
rect 10447 14692 10457 14703
rect 10457 14692 10503 14703
rect 10589 14692 10645 14748
rect 10731 14703 10787 14748
rect 10873 14703 10929 14748
rect 11015 14703 11071 14748
rect 10731 14692 10777 14703
rect 10777 14692 10787 14703
rect 10873 14692 10901 14703
rect 10901 14692 10929 14703
rect 11015 14692 11025 14703
rect 11025 14692 11071 14703
rect 10163 14579 10219 14606
rect 10305 14579 10361 14606
rect 10447 14579 10503 14606
rect 10163 14550 10209 14579
rect 10209 14550 10219 14579
rect 10305 14550 10333 14579
rect 10333 14550 10361 14579
rect 10447 14550 10457 14579
rect 10457 14550 10503 14579
rect 10589 14550 10645 14606
rect 10731 14579 10787 14606
rect 10873 14579 10929 14606
rect 11015 14579 11071 14606
rect 10731 14550 10777 14579
rect 10777 14550 10787 14579
rect 10873 14550 10901 14579
rect 10901 14550 10929 14579
rect 11015 14550 11025 14579
rect 11025 14550 11071 14579
rect 10163 14455 10219 14464
rect 10305 14455 10361 14464
rect 10447 14455 10503 14464
rect 10163 14408 10209 14455
rect 10209 14408 10219 14455
rect 10305 14408 10333 14455
rect 10333 14408 10361 14455
rect 10447 14408 10457 14455
rect 10457 14408 10503 14455
rect 10589 14408 10645 14464
rect 10731 14455 10787 14464
rect 10873 14455 10929 14464
rect 11015 14455 11071 14464
rect 10731 14408 10777 14455
rect 10777 14408 10787 14455
rect 10873 14408 10901 14455
rect 10901 14408 10929 14455
rect 11015 14408 11025 14455
rect 11025 14408 11071 14455
rect 11575 14699 11631 14755
rect 11717 14699 11773 14755
rect 11859 14699 11915 14755
rect 11575 14557 11631 14613
rect 11717 14557 11773 14613
rect 11859 14557 11915 14613
rect 11575 14415 11631 14471
rect 11717 14415 11773 14471
rect 11859 14415 11915 14471
rect 446 14273 502 14329
rect 588 14273 644 14329
rect 730 14273 786 14329
rect 446 14131 502 14187
rect 588 14131 644 14187
rect 730 14131 786 14187
rect 446 13989 502 14045
rect 588 13989 644 14045
rect 730 13989 786 14045
rect 446 13847 502 13903
rect 588 13847 644 13903
rect 730 13847 786 13903
rect 446 13705 502 13761
rect 588 13705 644 13761
rect 730 13705 786 13761
rect 446 13563 502 13619
rect 588 13563 644 13619
rect 730 13563 786 13619
rect 446 13421 502 13477
rect 588 13421 644 13477
rect 730 13421 786 13477
rect 11575 14273 11631 14329
rect 11717 14273 11773 14329
rect 11859 14273 11915 14329
rect 11575 14131 11631 14187
rect 11717 14131 11773 14187
rect 11859 14131 11915 14187
rect 11575 13989 11631 14045
rect 11717 13989 11773 14045
rect 11859 13989 11915 14045
rect 11575 13847 11631 13903
rect 11717 13847 11773 13903
rect 11859 13847 11915 13903
rect 11575 13705 11631 13761
rect 11717 13705 11773 13761
rect 11859 13705 11915 13761
rect 11575 13563 11631 13619
rect 11717 13563 11773 13619
rect 11859 13563 11915 13619
rect 11575 13421 11631 13477
rect 11717 13421 11773 13477
rect 11859 13421 11915 13477
rect 452 13109 508 13148
rect 594 13109 650 13148
rect 736 13109 792 13148
rect 452 13092 472 13109
rect 472 13092 508 13109
rect 594 13092 596 13109
rect 596 13092 648 13109
rect 648 13092 650 13109
rect 736 13092 772 13109
rect 772 13092 792 13109
rect 452 12985 508 13006
rect 594 12985 650 13006
rect 736 12985 792 13006
rect 452 12950 472 12985
rect 472 12950 508 12985
rect 594 12950 596 12985
rect 596 12950 648 12985
rect 648 12950 650 12985
rect 736 12950 772 12985
rect 772 12950 792 12985
rect 452 12861 508 12864
rect 594 12861 650 12864
rect 736 12861 792 12864
rect 452 12809 472 12861
rect 472 12809 508 12861
rect 594 12809 596 12861
rect 596 12809 648 12861
rect 648 12809 650 12861
rect 736 12809 772 12861
rect 772 12809 792 12861
rect 452 12808 508 12809
rect 594 12808 650 12809
rect 736 12808 792 12809
rect 452 12685 472 12722
rect 472 12685 508 12722
rect 594 12685 596 12722
rect 596 12685 648 12722
rect 648 12685 650 12722
rect 736 12685 772 12722
rect 772 12685 792 12722
rect 452 12666 508 12685
rect 594 12666 650 12685
rect 736 12666 792 12685
rect 452 12561 472 12580
rect 472 12561 508 12580
rect 594 12561 596 12580
rect 596 12561 648 12580
rect 648 12561 650 12580
rect 736 12561 772 12580
rect 772 12561 792 12580
rect 452 12524 508 12561
rect 594 12524 650 12561
rect 736 12524 792 12561
rect 452 12437 472 12438
rect 472 12437 508 12438
rect 594 12437 596 12438
rect 596 12437 648 12438
rect 648 12437 650 12438
rect 736 12437 772 12438
rect 772 12437 792 12438
rect 452 12382 508 12437
rect 594 12382 650 12437
rect 736 12382 792 12437
rect 452 12241 508 12296
rect 594 12241 650 12296
rect 736 12241 792 12296
rect 452 12240 472 12241
rect 472 12240 508 12241
rect 594 12240 596 12241
rect 596 12240 648 12241
rect 648 12240 650 12241
rect 736 12240 772 12241
rect 772 12240 792 12241
rect 452 12117 508 12154
rect 594 12117 650 12154
rect 736 12117 792 12154
rect 452 12098 472 12117
rect 472 12098 508 12117
rect 594 12098 596 12117
rect 596 12098 648 12117
rect 648 12098 650 12117
rect 736 12098 772 12117
rect 772 12098 792 12117
rect 452 11993 508 12012
rect 594 11993 650 12012
rect 736 11993 792 12012
rect 452 11956 472 11993
rect 472 11956 508 11993
rect 594 11956 596 11993
rect 596 11956 648 11993
rect 648 11956 650 11993
rect 736 11956 772 11993
rect 772 11956 792 11993
rect 452 11869 508 11870
rect 594 11869 650 11870
rect 736 11869 792 11870
rect 452 11817 472 11869
rect 472 11817 508 11869
rect 594 11817 596 11869
rect 596 11817 648 11869
rect 648 11817 650 11869
rect 736 11817 772 11869
rect 772 11817 792 11869
rect 452 11814 508 11817
rect 594 11814 650 11817
rect 736 11814 792 11817
rect 452 11693 472 11728
rect 472 11693 508 11728
rect 594 11693 596 11728
rect 596 11693 648 11728
rect 648 11693 650 11728
rect 736 11693 772 11728
rect 772 11693 792 11728
rect 452 11672 508 11693
rect 594 11672 650 11693
rect 736 11672 792 11693
rect 452 11569 472 11586
rect 472 11569 508 11586
rect 594 11569 596 11586
rect 596 11569 648 11586
rect 648 11569 650 11586
rect 736 11569 772 11586
rect 772 11569 792 11586
rect 452 11530 508 11569
rect 594 11530 650 11569
rect 736 11530 792 11569
rect 11581 13109 11637 13148
rect 11723 13109 11779 13148
rect 11865 13109 11921 13148
rect 11581 13092 11601 13109
rect 11601 13092 11637 13109
rect 11723 13092 11725 13109
rect 11725 13092 11777 13109
rect 11777 13092 11779 13109
rect 11865 13092 11901 13109
rect 11901 13092 11921 13109
rect 11581 12985 11637 13006
rect 11723 12985 11779 13006
rect 11865 12985 11921 13006
rect 11581 12950 11601 12985
rect 11601 12950 11637 12985
rect 11723 12950 11725 12985
rect 11725 12950 11777 12985
rect 11777 12950 11779 12985
rect 11865 12950 11901 12985
rect 11901 12950 11921 12985
rect 11581 12861 11637 12864
rect 11723 12861 11779 12864
rect 11865 12861 11921 12864
rect 11581 12809 11601 12861
rect 11601 12809 11637 12861
rect 11723 12809 11725 12861
rect 11725 12809 11777 12861
rect 11777 12809 11779 12861
rect 11865 12809 11901 12861
rect 11901 12809 11921 12861
rect 11581 12808 11637 12809
rect 11723 12808 11779 12809
rect 11865 12808 11921 12809
rect 11581 12685 11601 12722
rect 11601 12685 11637 12722
rect 11723 12685 11725 12722
rect 11725 12685 11777 12722
rect 11777 12685 11779 12722
rect 11865 12685 11901 12722
rect 11901 12685 11921 12722
rect 11581 12666 11637 12685
rect 11723 12666 11779 12685
rect 11865 12666 11921 12685
rect 11581 12561 11601 12580
rect 11601 12561 11637 12580
rect 11723 12561 11725 12580
rect 11725 12561 11777 12580
rect 11777 12561 11779 12580
rect 11865 12561 11901 12580
rect 11901 12561 11921 12580
rect 11581 12524 11637 12561
rect 11723 12524 11779 12561
rect 11865 12524 11921 12561
rect 11581 12437 11601 12438
rect 11601 12437 11637 12438
rect 11723 12437 11725 12438
rect 11725 12437 11777 12438
rect 11777 12437 11779 12438
rect 11865 12437 11901 12438
rect 11901 12437 11921 12438
rect 11581 12382 11637 12437
rect 11723 12382 11779 12437
rect 11865 12382 11921 12437
rect 11581 12241 11637 12296
rect 11723 12241 11779 12296
rect 11865 12241 11921 12296
rect 11581 12240 11601 12241
rect 11601 12240 11637 12241
rect 11723 12240 11725 12241
rect 11725 12240 11777 12241
rect 11777 12240 11779 12241
rect 11865 12240 11901 12241
rect 11901 12240 11921 12241
rect 11581 12117 11637 12154
rect 11723 12117 11779 12154
rect 11865 12117 11921 12154
rect 11581 12098 11601 12117
rect 11601 12098 11637 12117
rect 11723 12098 11725 12117
rect 11725 12098 11777 12117
rect 11777 12098 11779 12117
rect 11865 12098 11901 12117
rect 11901 12098 11921 12117
rect 11581 11993 11637 12012
rect 11723 11993 11779 12012
rect 11865 11993 11921 12012
rect 11581 11956 11601 11993
rect 11601 11956 11637 11993
rect 11723 11956 11725 11993
rect 11725 11956 11777 11993
rect 11777 11956 11779 11993
rect 11865 11956 11901 11993
rect 11901 11956 11921 11993
rect 11581 11869 11637 11870
rect 11723 11869 11779 11870
rect 11865 11869 11921 11870
rect 11581 11817 11601 11869
rect 11601 11817 11637 11869
rect 11723 11817 11725 11869
rect 11725 11817 11777 11869
rect 11777 11817 11779 11869
rect 11865 11817 11901 11869
rect 11901 11817 11921 11869
rect 11581 11814 11637 11817
rect 11723 11814 11779 11817
rect 11865 11814 11921 11817
rect 11581 11693 11601 11728
rect 11601 11693 11637 11728
rect 11723 11693 11725 11728
rect 11725 11693 11777 11728
rect 11777 11693 11779 11728
rect 11865 11693 11901 11728
rect 11901 11693 11921 11728
rect 11581 11672 11637 11693
rect 11723 11672 11779 11693
rect 11865 11672 11921 11693
rect 11581 11569 11601 11586
rect 11601 11569 11637 11586
rect 11723 11569 11725 11586
rect 11725 11569 11777 11586
rect 11777 11569 11779 11586
rect 11865 11569 11901 11586
rect 11901 11569 11921 11586
rect 11581 11530 11637 11569
rect 11723 11530 11779 11569
rect 11865 11530 11921 11569
rect 471 10861 527 10887
rect 613 10861 669 10887
rect 471 10831 527 10861
rect 613 10831 669 10861
rect 471 10689 527 10745
rect 613 10689 669 10745
rect 471 10547 527 10603
rect 613 10547 669 10603
rect 471 10405 527 10461
rect 613 10405 669 10461
rect 471 10289 527 10319
rect 613 10289 669 10319
rect 471 10263 527 10289
rect 613 10263 669 10289
rect 11713 10861 11769 10887
rect 11855 10861 11911 10887
rect 11713 10831 11769 10861
rect 11855 10831 11911 10861
rect 11713 10689 11769 10745
rect 11855 10689 11911 10745
rect 11713 10547 11769 10603
rect 11855 10547 11911 10603
rect 11713 10405 11769 10461
rect 11855 10405 11911 10461
rect 11713 10289 11769 10319
rect 11855 10289 11911 10319
rect 11713 10263 11769 10289
rect 11855 10263 11911 10289
rect 471 9866 527 9922
rect 613 9866 669 9922
rect 471 9724 527 9780
rect 613 9724 669 9780
rect 471 9582 527 9638
rect 613 9582 669 9638
rect 471 9440 527 9496
rect 613 9440 669 9496
rect 471 9298 527 9354
rect 613 9298 669 9354
rect 471 9156 527 9212
rect 613 9156 669 9212
rect 471 9014 527 9070
rect 613 9014 669 9070
rect 471 8872 527 8928
rect 613 8872 669 8928
rect 471 8730 527 8786
rect 613 8730 669 8786
rect 471 8588 527 8644
rect 613 8588 669 8644
rect 471 8446 527 8502
rect 613 8446 669 8502
rect 471 8304 527 8360
rect 613 8304 669 8360
rect 471 8162 527 8218
rect 613 8162 669 8218
rect 471 8020 527 8076
rect 613 8020 669 8076
rect 471 7878 527 7934
rect 613 7878 669 7934
rect 471 7736 527 7792
rect 613 7736 669 7792
rect 471 7594 527 7650
rect 613 7594 669 7650
rect 471 7452 527 7508
rect 613 7452 669 7508
rect 471 7310 527 7366
rect 613 7310 669 7366
rect 471 7168 527 7224
rect 613 7168 669 7224
rect 471 7026 527 7082
rect 613 7026 669 7082
rect 11713 9866 11769 9922
rect 11855 9866 11911 9922
rect 11713 9724 11769 9780
rect 11855 9724 11911 9780
rect 11713 9582 11769 9638
rect 11855 9582 11911 9638
rect 11713 9440 11769 9496
rect 11855 9440 11911 9496
rect 11713 9298 11769 9354
rect 11855 9298 11911 9354
rect 11713 9156 11769 9212
rect 11855 9156 11911 9212
rect 11713 9014 11769 9070
rect 11855 9014 11911 9070
rect 11713 8872 11769 8928
rect 11855 8872 11911 8928
rect 11713 8730 11769 8786
rect 11855 8730 11911 8786
rect 11713 8588 11769 8644
rect 11855 8588 11911 8644
rect 11713 8446 11769 8502
rect 11855 8446 11911 8502
rect 11713 8304 11769 8360
rect 11855 8304 11911 8360
rect 11713 8162 11769 8218
rect 11855 8162 11911 8218
rect 11713 8020 11769 8076
rect 11855 8020 11911 8076
rect 11713 7878 11769 7934
rect 11855 7878 11911 7934
rect 11713 7736 11769 7792
rect 11855 7736 11911 7792
rect 11713 7594 11769 7650
rect 11855 7594 11911 7650
rect 11713 7452 11769 7508
rect 11855 7452 11911 7508
rect 11713 7310 11769 7366
rect 11855 7310 11911 7366
rect 11713 7168 11769 7224
rect 11855 7168 11911 7224
rect 11713 7026 11769 7082
rect 11855 7026 11911 7082
rect 471 6684 527 6740
rect 613 6684 669 6740
rect 471 6542 527 6598
rect 613 6542 669 6598
rect 471 6400 527 6456
rect 613 6400 669 6456
rect 471 6258 527 6314
rect 613 6258 669 6314
rect 471 6116 527 6172
rect 613 6116 669 6172
rect 471 5974 527 6030
rect 613 5974 669 6030
rect 471 5832 527 5888
rect 613 5832 669 5888
rect 471 5690 527 5746
rect 613 5690 669 5746
rect 471 5548 527 5604
rect 613 5548 669 5604
rect 471 5406 527 5462
rect 613 5406 669 5462
rect 471 5264 527 5320
rect 613 5264 669 5320
rect 471 5122 527 5178
rect 613 5122 669 5178
rect 471 4980 527 5036
rect 613 4980 669 5036
rect 471 4838 527 4894
rect 613 4838 669 4894
rect 471 4696 527 4752
rect 613 4696 669 4752
rect 471 4554 527 4610
rect 613 4554 669 4610
rect 471 4412 527 4468
rect 613 4412 669 4468
rect 471 4270 527 4326
rect 613 4270 669 4326
rect 471 4128 527 4184
rect 613 4128 669 4184
rect 471 3986 527 4042
rect 613 3986 669 4042
rect 471 3844 527 3900
rect 613 3844 669 3900
rect 11713 6684 11769 6740
rect 11855 6684 11911 6740
rect 11713 6542 11769 6598
rect 11855 6542 11911 6598
rect 11713 6400 11769 6456
rect 11855 6400 11911 6456
rect 11713 6258 11769 6314
rect 11855 6258 11911 6314
rect 11713 6116 11769 6172
rect 11855 6116 11911 6172
rect 11713 5974 11769 6030
rect 11855 5974 11911 6030
rect 11713 5832 11769 5888
rect 11855 5832 11911 5888
rect 11713 5690 11769 5746
rect 11855 5690 11911 5746
rect 11713 5548 11769 5604
rect 11855 5548 11911 5604
rect 11713 5406 11769 5462
rect 11855 5406 11911 5462
rect 11713 5264 11769 5320
rect 11855 5264 11911 5320
rect 11713 5122 11769 5178
rect 11855 5122 11911 5178
rect 11713 4980 11769 5036
rect 11855 4980 11911 5036
rect 11713 4838 11769 4894
rect 11855 4838 11911 4894
rect 11713 4696 11769 4752
rect 11855 4696 11911 4752
rect 11713 4554 11769 4610
rect 11855 4554 11911 4610
rect 11713 4412 11769 4468
rect 11855 4412 11911 4468
rect 11713 4270 11769 4326
rect 11855 4270 11911 4326
rect 11713 4128 11769 4184
rect 11855 4128 11911 4184
rect 11713 3986 11769 4042
rect 11855 3986 11911 4042
rect 11713 3844 11769 3900
rect 11855 3844 11911 3900
rect 471 3505 527 3522
rect 613 3505 669 3522
rect 471 3466 527 3505
rect 613 3466 669 3505
rect 471 3324 527 3380
rect 613 3324 669 3380
rect 471 3182 527 3238
rect 613 3182 669 3238
rect 471 3040 527 3096
rect 613 3040 669 3096
rect 11713 3505 11769 3522
rect 11855 3505 11911 3522
rect 11713 3466 11769 3505
rect 11855 3466 11911 3505
rect 11713 3324 11769 3380
rect 11855 3324 11911 3380
rect 11713 3182 11769 3238
rect 11855 3182 11911 3238
rect 11713 3040 11769 3096
rect 11855 3040 11911 3096
rect 452 2278 508 2317
rect 594 2278 650 2317
rect 736 2278 792 2317
rect 452 2261 472 2278
rect 472 2261 508 2278
rect 594 2261 596 2278
rect 596 2261 648 2278
rect 648 2261 650 2278
rect 736 2261 772 2278
rect 772 2261 792 2278
rect 452 2154 508 2175
rect 594 2154 650 2175
rect 736 2154 792 2175
rect 452 2119 472 2154
rect 472 2119 508 2154
rect 594 2119 596 2154
rect 596 2119 648 2154
rect 648 2119 650 2154
rect 736 2119 772 2154
rect 772 2119 792 2154
rect 452 2030 508 2033
rect 594 2030 650 2033
rect 736 2030 792 2033
rect 452 1978 472 2030
rect 472 1978 508 2030
rect 594 1978 596 2030
rect 596 1978 648 2030
rect 648 1978 650 2030
rect 736 1978 772 2030
rect 772 1978 792 2030
rect 452 1977 508 1978
rect 594 1977 650 1978
rect 736 1977 792 1978
rect 452 1854 472 1891
rect 472 1854 508 1891
rect 594 1854 596 1891
rect 596 1854 648 1891
rect 648 1854 650 1891
rect 736 1854 772 1891
rect 772 1854 792 1891
rect 452 1835 508 1854
rect 594 1835 650 1854
rect 736 1835 792 1854
rect 452 1730 472 1749
rect 472 1730 508 1749
rect 594 1730 596 1749
rect 596 1730 648 1749
rect 648 1730 650 1749
rect 736 1730 772 1749
rect 772 1730 792 1749
rect 452 1693 508 1730
rect 594 1693 650 1730
rect 736 1693 792 1730
rect 452 1606 472 1607
rect 472 1606 508 1607
rect 594 1606 596 1607
rect 596 1606 648 1607
rect 648 1606 650 1607
rect 736 1606 772 1607
rect 772 1606 792 1607
rect 452 1551 508 1606
rect 594 1551 650 1606
rect 736 1551 792 1606
rect 452 1410 508 1465
rect 594 1410 650 1465
rect 736 1410 792 1465
rect 452 1409 472 1410
rect 472 1409 508 1410
rect 594 1409 596 1410
rect 596 1409 648 1410
rect 648 1409 650 1410
rect 736 1409 772 1410
rect 772 1409 792 1410
rect 452 1286 508 1323
rect 594 1286 650 1323
rect 736 1286 792 1323
rect 452 1267 472 1286
rect 472 1267 508 1286
rect 594 1267 596 1286
rect 596 1267 648 1286
rect 648 1267 650 1286
rect 736 1267 772 1286
rect 772 1267 792 1286
rect 452 1162 508 1181
rect 594 1162 650 1181
rect 736 1162 792 1181
rect 452 1125 472 1162
rect 472 1125 508 1162
rect 594 1125 596 1162
rect 596 1125 648 1162
rect 648 1125 650 1162
rect 736 1125 772 1162
rect 772 1125 792 1162
rect 452 1038 508 1039
rect 594 1038 650 1039
rect 736 1038 792 1039
rect 452 986 472 1038
rect 472 986 508 1038
rect 594 986 596 1038
rect 596 986 648 1038
rect 648 986 650 1038
rect 736 986 772 1038
rect 772 986 792 1038
rect 452 983 508 986
rect 594 983 650 986
rect 736 983 792 986
rect 452 862 472 897
rect 472 862 508 897
rect 594 862 596 897
rect 596 862 648 897
rect 648 862 650 897
rect 736 862 772 897
rect 772 862 792 897
rect 452 841 508 862
rect 594 841 650 862
rect 736 841 792 862
rect 452 738 472 755
rect 472 738 508 755
rect 594 738 596 755
rect 596 738 648 755
rect 648 738 650 755
rect 736 738 772 755
rect 772 738 792 755
rect 452 699 508 738
rect 594 699 650 738
rect 736 699 792 738
rect 11581 2278 11637 2317
rect 11723 2278 11779 2317
rect 11865 2278 11921 2317
rect 11581 2261 11601 2278
rect 11601 2261 11637 2278
rect 11723 2261 11725 2278
rect 11725 2261 11777 2278
rect 11777 2261 11779 2278
rect 11865 2261 11901 2278
rect 11901 2261 11921 2278
rect 11581 2154 11637 2175
rect 11723 2154 11779 2175
rect 11865 2154 11921 2175
rect 11581 2119 11601 2154
rect 11601 2119 11637 2154
rect 11723 2119 11725 2154
rect 11725 2119 11777 2154
rect 11777 2119 11779 2154
rect 11865 2119 11901 2154
rect 11901 2119 11921 2154
rect 11581 2030 11637 2033
rect 11723 2030 11779 2033
rect 11865 2030 11921 2033
rect 11581 1978 11601 2030
rect 11601 1978 11637 2030
rect 11723 1978 11725 2030
rect 11725 1978 11777 2030
rect 11777 1978 11779 2030
rect 11865 1978 11901 2030
rect 11901 1978 11921 2030
rect 11581 1977 11637 1978
rect 11723 1977 11779 1978
rect 11865 1977 11921 1978
rect 11581 1854 11601 1891
rect 11601 1854 11637 1891
rect 11723 1854 11725 1891
rect 11725 1854 11777 1891
rect 11777 1854 11779 1891
rect 11865 1854 11901 1891
rect 11901 1854 11921 1891
rect 11581 1835 11637 1854
rect 11723 1835 11779 1854
rect 11865 1835 11921 1854
rect 11581 1730 11601 1749
rect 11601 1730 11637 1749
rect 11723 1730 11725 1749
rect 11725 1730 11777 1749
rect 11777 1730 11779 1749
rect 11865 1730 11901 1749
rect 11901 1730 11921 1749
rect 11581 1693 11637 1730
rect 11723 1693 11779 1730
rect 11865 1693 11921 1730
rect 11581 1606 11601 1607
rect 11601 1606 11637 1607
rect 11723 1606 11725 1607
rect 11725 1606 11777 1607
rect 11777 1606 11779 1607
rect 11865 1606 11901 1607
rect 11901 1606 11921 1607
rect 11581 1551 11637 1606
rect 11723 1551 11779 1606
rect 11865 1551 11921 1606
rect 11581 1410 11637 1465
rect 11723 1410 11779 1465
rect 11865 1410 11921 1465
rect 11581 1409 11601 1410
rect 11601 1409 11637 1410
rect 11723 1409 11725 1410
rect 11725 1409 11777 1410
rect 11777 1409 11779 1410
rect 11865 1409 11901 1410
rect 11901 1409 11921 1410
rect 11581 1286 11637 1323
rect 11723 1286 11779 1323
rect 11865 1286 11921 1323
rect 11581 1267 11601 1286
rect 11601 1267 11637 1286
rect 11723 1267 11725 1286
rect 11725 1267 11777 1286
rect 11777 1267 11779 1286
rect 11865 1267 11901 1286
rect 11901 1267 11921 1286
rect 11581 1162 11637 1181
rect 11723 1162 11779 1181
rect 11865 1162 11921 1181
rect 11581 1125 11601 1162
rect 11601 1125 11637 1162
rect 11723 1125 11725 1162
rect 11725 1125 11777 1162
rect 11777 1125 11779 1162
rect 11865 1125 11901 1162
rect 11901 1125 11921 1162
rect 11581 1038 11637 1039
rect 11723 1038 11779 1039
rect 11865 1038 11921 1039
rect 11581 986 11601 1038
rect 11601 986 11637 1038
rect 11723 986 11725 1038
rect 11725 986 11777 1038
rect 11777 986 11779 1038
rect 11865 986 11901 1038
rect 11901 986 11921 1038
rect 11581 983 11637 986
rect 11723 983 11779 986
rect 11865 983 11921 986
rect 11581 862 11601 897
rect 11601 862 11637 897
rect 11723 862 11725 897
rect 11725 862 11777 897
rect 11777 862 11779 897
rect 11865 862 11901 897
rect 11901 862 11921 897
rect 11581 841 11637 862
rect 11723 841 11779 862
rect 11865 841 11921 862
rect 11581 738 11601 755
rect 11601 738 11637 755
rect 11723 738 11725 755
rect 11725 738 11777 755
rect 11777 738 11779 755
rect 11865 738 11901 755
rect 11901 738 11921 755
rect 11581 699 11637 738
rect 11723 699 11779 738
rect 11865 699 11921 738
rect 12870 339 12926 356
rect 13012 339 13068 356
rect 12870 300 12891 339
rect 12891 300 12926 339
rect 13012 300 13047 339
rect 13047 300 13068 339
rect -717 232 -696 288
rect -696 232 -661 288
rect -575 232 -540 288
rect -540 232 -519 288
rect -717 90 -696 146
rect -696 90 -661 146
rect -575 90 -540 146
rect -540 90 -519 146
rect -717 -52 -696 4
rect -696 -52 -661 4
rect -575 -52 -540 4
rect -540 -52 -519 4
rect -717 -194 -696 -138
rect -696 -194 -661 -138
rect -575 -194 -540 -138
rect -540 -194 -519 -138
rect -717 -336 -696 -280
rect -696 -336 -661 -280
rect -575 -336 -540 -280
rect -540 -336 -519 -280
rect -717 -478 -696 -422
rect -696 -478 -661 -422
rect -575 -478 -540 -422
rect -540 -478 -519 -422
rect -717 -620 -696 -564
rect -696 -620 -661 -564
rect -575 -620 -540 -564
rect -540 -620 -519 -564
rect -717 -762 -696 -706
rect -696 -762 -661 -706
rect -575 -762 -540 -706
rect -540 -762 -519 -706
rect -717 -904 -696 -848
rect -696 -904 -661 -848
rect -575 -904 -540 -848
rect -540 -904 -519 -848
rect 12870 158 12891 214
rect 12891 158 12926 214
rect 13012 158 13047 214
rect 13047 158 13068 214
rect 12870 16 12891 72
rect 12891 16 12926 72
rect 13012 16 13047 72
rect 13047 16 13068 72
rect 12870 -126 12891 -70
rect 12891 -126 12926 -70
rect 13012 -126 13047 -70
rect 13047 -126 13068 -70
rect 12870 -268 12891 -212
rect 12891 -268 12926 -212
rect 13012 -268 13047 -212
rect 13047 -268 13068 -212
rect 12870 -410 12891 -354
rect 12891 -410 12926 -354
rect 13012 -410 13047 -354
rect 13047 -410 13068 -354
rect 12870 -552 12891 -496
rect 12891 -552 12926 -496
rect 13012 -552 13047 -496
rect 13047 -552 13068 -496
rect 12870 -694 12891 -638
rect 12891 -694 12926 -638
rect 13012 -694 13047 -638
rect 13047 -694 13068 -638
rect 12870 -836 12891 -780
rect 12891 -836 12926 -780
rect 13012 -836 13047 -780
rect 13047 -836 13068 -780
rect 12870 -961 12891 -922
rect 12891 -961 12926 -922
rect 13012 -961 13047 -922
rect 13047 -961 13068 -922
rect 12870 -978 12926 -961
rect 13012 -978 13068 -961
<< metal3 >>
rect -694 14755 -476 14765
rect -694 14699 -684 14755
rect -628 14699 -542 14755
rect -486 14699 -476 14755
rect -694 14613 -476 14699
rect -694 14557 -684 14613
rect -628 14557 -542 14613
rect -486 14557 -476 14613
rect -694 14471 -476 14557
rect -694 14415 -684 14471
rect -628 14415 -542 14471
rect -486 14415 -476 14471
rect -694 14329 -476 14415
rect -694 14273 -684 14329
rect -628 14273 -542 14329
rect -486 14273 -476 14329
rect -694 14187 -476 14273
rect -694 14131 -684 14187
rect -628 14131 -542 14187
rect -486 14131 -476 14187
rect -694 14045 -476 14131
rect -694 13989 -684 14045
rect -628 13989 -542 14045
rect -486 13989 -476 14045
rect -694 13903 -476 13989
rect -694 13847 -684 13903
rect -628 13847 -542 13903
rect -486 13847 -476 13903
rect -694 13761 -476 13847
rect -694 13705 -684 13761
rect -628 13705 -542 13761
rect -486 13705 -476 13761
rect -694 13619 -476 13705
rect -694 13563 -684 13619
rect -628 13563 -542 13619
rect -486 13563 -476 13619
rect -694 13477 -476 13563
rect -694 13421 -684 13477
rect -628 13421 -542 13477
rect -486 13421 -476 13477
rect -694 13411 -476 13421
rect 436 14755 796 14765
rect 436 14699 446 14755
rect 502 14699 588 14755
rect 644 14699 730 14755
rect 786 14699 796 14755
rect 436 14613 796 14699
rect 436 14557 446 14613
rect 502 14557 588 14613
rect 644 14557 730 14613
rect 786 14557 796 14613
rect 436 14471 796 14557
rect 436 14415 446 14471
rect 502 14415 588 14471
rect 644 14415 730 14471
rect 786 14415 796 14471
rect 436 14329 796 14415
rect 1312 14748 2240 14758
rect 1312 14692 1322 14748
rect 1378 14692 1464 14748
rect 1520 14692 1606 14748
rect 1662 14692 1748 14748
rect 1804 14692 1890 14748
rect 1946 14692 2032 14748
rect 2088 14692 2174 14748
rect 2230 14692 2240 14748
rect 1312 14606 2240 14692
rect 1312 14550 1322 14606
rect 1378 14550 1464 14606
rect 1520 14550 1606 14606
rect 1662 14550 1748 14606
rect 1804 14550 1890 14606
rect 1946 14550 2032 14606
rect 2088 14550 2174 14606
rect 2230 14550 2240 14606
rect 1312 14464 2240 14550
rect 1312 14408 1322 14464
rect 1378 14408 1464 14464
rect 1520 14408 1606 14464
rect 1662 14408 1748 14464
rect 1804 14408 1890 14464
rect 1946 14408 2032 14464
rect 2088 14408 2174 14464
rect 2230 14408 2240 14464
rect 1312 14398 2240 14408
rect 3084 14748 4012 14758
rect 3084 14692 3094 14748
rect 3150 14692 3236 14748
rect 3292 14692 3378 14748
rect 3434 14692 3520 14748
rect 3576 14692 3662 14748
rect 3718 14692 3804 14748
rect 3860 14692 3946 14748
rect 4002 14692 4012 14748
rect 3084 14606 4012 14692
rect 3084 14550 3094 14606
rect 3150 14550 3236 14606
rect 3292 14550 3378 14606
rect 3434 14550 3520 14606
rect 3576 14550 3662 14606
rect 3718 14550 3804 14606
rect 3860 14550 3946 14606
rect 4002 14550 4012 14606
rect 3084 14464 4012 14550
rect 3084 14408 3094 14464
rect 3150 14408 3236 14464
rect 3292 14408 3378 14464
rect 3434 14408 3520 14464
rect 3576 14408 3662 14464
rect 3718 14408 3804 14464
rect 3860 14408 3946 14464
rect 4002 14408 4012 14464
rect 3084 14398 4012 14408
rect 4849 14748 5777 14758
rect 4849 14692 4859 14748
rect 4915 14692 5001 14748
rect 5057 14692 5143 14748
rect 5199 14692 5285 14748
rect 5341 14692 5427 14748
rect 5483 14692 5569 14748
rect 5625 14692 5711 14748
rect 5767 14692 5777 14748
rect 4849 14606 5777 14692
rect 4849 14550 4859 14606
rect 4915 14550 5001 14606
rect 5057 14550 5143 14606
rect 5199 14550 5285 14606
rect 5341 14550 5427 14606
rect 5483 14550 5569 14606
rect 5625 14550 5711 14606
rect 5767 14550 5777 14606
rect 4849 14464 5777 14550
rect 4849 14408 4859 14464
rect 4915 14408 5001 14464
rect 5057 14408 5143 14464
rect 5199 14408 5285 14464
rect 5341 14408 5427 14464
rect 5483 14408 5569 14464
rect 5625 14408 5711 14464
rect 5767 14408 5777 14464
rect 4849 14398 5777 14408
rect 6618 14748 7546 14758
rect 6618 14692 6628 14748
rect 6684 14692 6770 14748
rect 6826 14692 6912 14748
rect 6968 14692 7054 14748
rect 7110 14692 7196 14748
rect 7252 14692 7338 14748
rect 7394 14692 7480 14748
rect 7536 14692 7546 14748
rect 6618 14606 7546 14692
rect 6618 14550 6628 14606
rect 6684 14550 6770 14606
rect 6826 14550 6912 14606
rect 6968 14550 7054 14606
rect 7110 14550 7196 14606
rect 7252 14550 7338 14606
rect 7394 14550 7480 14606
rect 7536 14550 7546 14606
rect 6618 14464 7546 14550
rect 6618 14408 6628 14464
rect 6684 14408 6770 14464
rect 6826 14408 6912 14464
rect 6968 14408 7054 14464
rect 7110 14408 7196 14464
rect 7252 14408 7338 14464
rect 7394 14408 7480 14464
rect 7536 14408 7546 14464
rect 6618 14398 7546 14408
rect 8387 14748 9315 14758
rect 8387 14692 8397 14748
rect 8453 14692 8539 14748
rect 8595 14692 8681 14748
rect 8737 14692 8823 14748
rect 8879 14692 8965 14748
rect 9021 14692 9107 14748
rect 9163 14692 9249 14748
rect 9305 14692 9315 14748
rect 8387 14606 9315 14692
rect 8387 14550 8397 14606
rect 8453 14550 8539 14606
rect 8595 14550 8681 14606
rect 8737 14550 8823 14606
rect 8879 14550 8965 14606
rect 9021 14550 9107 14606
rect 9163 14550 9249 14606
rect 9305 14550 9315 14606
rect 8387 14464 9315 14550
rect 8387 14408 8397 14464
rect 8453 14408 8539 14464
rect 8595 14408 8681 14464
rect 8737 14408 8823 14464
rect 8879 14408 8965 14464
rect 9021 14408 9107 14464
rect 9163 14408 9249 14464
rect 9305 14408 9315 14464
rect 8387 14398 9315 14408
rect 10153 14748 11081 14758
rect 10153 14692 10163 14748
rect 10219 14692 10305 14748
rect 10361 14692 10447 14748
rect 10503 14692 10589 14748
rect 10645 14692 10731 14748
rect 10787 14692 10873 14748
rect 10929 14692 11015 14748
rect 11071 14692 11081 14748
rect 10153 14606 11081 14692
rect 10153 14550 10163 14606
rect 10219 14550 10305 14606
rect 10361 14550 10447 14606
rect 10503 14550 10589 14606
rect 10645 14550 10731 14606
rect 10787 14550 10873 14606
rect 10929 14550 11015 14606
rect 11071 14550 11081 14606
rect 10153 14464 11081 14550
rect 10153 14408 10163 14464
rect 10219 14408 10305 14464
rect 10361 14408 10447 14464
rect 10503 14408 10589 14464
rect 10645 14408 10731 14464
rect 10787 14408 10873 14464
rect 10929 14408 11015 14464
rect 11071 14408 11081 14464
rect 10153 14398 11081 14408
rect 11565 14755 11925 14765
rect 11565 14699 11575 14755
rect 11631 14699 11717 14755
rect 11773 14699 11859 14755
rect 11915 14699 11925 14755
rect 11565 14613 11925 14699
rect 11565 14557 11575 14613
rect 11631 14557 11717 14613
rect 11773 14557 11859 14613
rect 11915 14557 11925 14613
rect 11565 14471 11925 14557
rect 11565 14415 11575 14471
rect 11631 14415 11717 14471
rect 11773 14415 11859 14471
rect 11915 14415 11925 14471
rect 436 14273 446 14329
rect 502 14273 588 14329
rect 644 14273 730 14329
rect 786 14273 796 14329
rect 436 14187 796 14273
rect 436 14131 446 14187
rect 502 14131 588 14187
rect 644 14131 730 14187
rect 786 14131 796 14187
rect 436 14045 796 14131
rect 436 13989 446 14045
rect 502 13989 588 14045
rect 644 13989 730 14045
rect 786 13989 796 14045
rect 436 13903 796 13989
rect 436 13847 446 13903
rect 502 13847 588 13903
rect 644 13847 730 13903
rect 786 13847 796 13903
rect 436 13761 796 13847
rect 436 13705 446 13761
rect 502 13705 588 13761
rect 644 13705 730 13761
rect 786 13705 796 13761
rect 436 13619 796 13705
rect 436 13563 446 13619
rect 502 13563 588 13619
rect 644 13563 730 13619
rect 786 13563 796 13619
rect 436 13477 796 13563
rect 436 13421 446 13477
rect 502 13421 588 13477
rect 644 13421 730 13477
rect 786 13421 796 13477
rect 436 13411 796 13421
rect 11565 14329 11925 14415
rect 11565 14273 11575 14329
rect 11631 14273 11717 14329
rect 11773 14273 11859 14329
rect 11915 14273 11925 14329
rect 11565 14187 11925 14273
rect 11565 14131 11575 14187
rect 11631 14131 11717 14187
rect 11773 14131 11859 14187
rect 11915 14131 11925 14187
rect 11565 14045 11925 14131
rect 11565 13989 11575 14045
rect 11631 13989 11717 14045
rect 11773 13989 11859 14045
rect 11915 13989 11925 14045
rect 11565 13903 11925 13989
rect 11565 13847 11575 13903
rect 11631 13847 11717 13903
rect 11773 13847 11859 13903
rect 11915 13847 11925 13903
rect 11565 13761 11925 13847
rect 11565 13705 11575 13761
rect 11631 13705 11717 13761
rect 11773 13705 11859 13761
rect 11915 13705 11925 13761
rect 11565 13619 11925 13705
rect 11565 13563 11575 13619
rect 11631 13563 11717 13619
rect 11773 13563 11859 13619
rect 11915 13563 11925 13619
rect 11565 13477 11925 13563
rect 11565 13421 11575 13477
rect 11631 13421 11717 13477
rect 11773 13421 11859 13477
rect 11915 13421 11925 13477
rect 11565 13411 11925 13421
rect 442 13148 802 13158
rect 442 13092 452 13148
rect 508 13092 594 13148
rect 650 13092 736 13148
rect 792 13092 802 13148
rect 442 13006 802 13092
rect 442 12950 452 13006
rect 508 12950 594 13006
rect 650 12950 736 13006
rect 792 12950 802 13006
rect 442 12864 802 12950
rect 442 12808 452 12864
rect 508 12808 594 12864
rect 650 12808 736 12864
rect 792 12808 802 12864
rect 442 12722 802 12808
rect 442 12666 452 12722
rect 508 12666 594 12722
rect 650 12666 736 12722
rect 792 12666 802 12722
rect 442 12580 802 12666
rect 442 12524 452 12580
rect 508 12524 594 12580
rect 650 12524 736 12580
rect 792 12524 802 12580
rect 442 12438 802 12524
rect 442 12382 452 12438
rect 508 12382 594 12438
rect 650 12382 736 12438
rect 792 12382 802 12438
rect 442 12296 802 12382
rect 442 12240 452 12296
rect 508 12240 594 12296
rect 650 12240 736 12296
rect 792 12240 802 12296
rect 442 12154 802 12240
rect 442 12098 452 12154
rect 508 12098 594 12154
rect 650 12098 736 12154
rect 792 12098 802 12154
rect 442 12012 802 12098
rect 442 11956 452 12012
rect 508 11956 594 12012
rect 650 11956 736 12012
rect 792 11956 802 12012
rect 442 11870 802 11956
rect 442 11814 452 11870
rect 508 11814 594 11870
rect 650 11814 736 11870
rect 792 11814 802 11870
rect 442 11728 802 11814
rect 442 11672 452 11728
rect 508 11672 594 11728
rect 650 11672 736 11728
rect 792 11672 802 11728
rect 442 11586 802 11672
rect 442 11530 452 11586
rect 508 11530 594 11586
rect 650 11530 736 11586
rect 792 11530 802 11586
rect 442 11520 802 11530
rect 11571 13148 11931 13158
rect 11571 13092 11581 13148
rect 11637 13092 11723 13148
rect 11779 13092 11865 13148
rect 11921 13092 11931 13148
rect 11571 13006 11931 13092
rect 11571 12950 11581 13006
rect 11637 12950 11723 13006
rect 11779 12950 11865 13006
rect 11921 12950 11931 13006
rect 11571 12864 11931 12950
rect 11571 12808 11581 12864
rect 11637 12808 11723 12864
rect 11779 12808 11865 12864
rect 11921 12808 11931 12864
rect 11571 12722 11931 12808
rect 11571 12666 11581 12722
rect 11637 12666 11723 12722
rect 11779 12666 11865 12722
rect 11921 12666 11931 12722
rect 11571 12580 11931 12666
rect 11571 12524 11581 12580
rect 11637 12524 11723 12580
rect 11779 12524 11865 12580
rect 11921 12524 11931 12580
rect 11571 12438 11931 12524
rect 11571 12382 11581 12438
rect 11637 12382 11723 12438
rect 11779 12382 11865 12438
rect 11921 12382 11931 12438
rect 11571 12296 11931 12382
rect 11571 12240 11581 12296
rect 11637 12240 11723 12296
rect 11779 12240 11865 12296
rect 11921 12240 11931 12296
rect 11571 12154 11931 12240
rect 11571 12098 11581 12154
rect 11637 12098 11723 12154
rect 11779 12098 11865 12154
rect 11921 12098 11931 12154
rect 11571 12012 11931 12098
rect 11571 11956 11581 12012
rect 11637 11956 11723 12012
rect 11779 11956 11865 12012
rect 11921 11956 11931 12012
rect 11571 11870 11931 11956
rect 11571 11814 11581 11870
rect 11637 11814 11723 11870
rect 11779 11814 11865 11870
rect 11921 11814 11931 11870
rect 11571 11728 11931 11814
rect 11571 11672 11581 11728
rect 11637 11672 11723 11728
rect 11779 11672 11865 11728
rect 11921 11672 11931 11728
rect 11571 11586 11931 11672
rect 11571 11530 11581 11586
rect 11637 11530 11723 11586
rect 11779 11530 11865 11586
rect 11921 11530 11931 11586
rect 11571 11520 11931 11530
rect 461 10887 679 10897
rect 461 10831 471 10887
rect 527 10831 613 10887
rect 669 10831 679 10887
rect 461 10745 679 10831
rect 461 10689 471 10745
rect 527 10689 613 10745
rect 669 10689 679 10745
rect 461 10603 679 10689
rect 461 10547 471 10603
rect 527 10547 613 10603
rect 669 10547 679 10603
rect 461 10461 679 10547
rect 461 10405 471 10461
rect 527 10405 613 10461
rect 669 10405 679 10461
rect 461 10319 679 10405
rect 461 10263 471 10319
rect 527 10263 613 10319
rect 669 10263 679 10319
rect 461 10253 679 10263
rect 11703 10887 11921 10897
rect 11703 10831 11713 10887
rect 11769 10831 11855 10887
rect 11911 10831 11921 10887
rect 11703 10745 11921 10831
rect 11703 10689 11713 10745
rect 11769 10689 11855 10745
rect 11911 10689 11921 10745
rect 11703 10603 11921 10689
rect 11703 10547 11713 10603
rect 11769 10547 11855 10603
rect 11911 10547 11921 10603
rect 11703 10461 11921 10547
rect 11703 10405 11713 10461
rect 11769 10405 11855 10461
rect 11911 10405 11921 10461
rect 11703 10319 11921 10405
rect 11703 10263 11713 10319
rect 11769 10263 11855 10319
rect 11911 10263 11921 10319
rect 11703 10253 11921 10263
rect 461 9922 679 9932
rect 461 9866 471 9922
rect 527 9866 613 9922
rect 669 9866 679 9922
rect 461 9780 679 9866
rect 461 9724 471 9780
rect 527 9724 613 9780
rect 669 9724 679 9780
rect 461 9638 679 9724
rect 461 9582 471 9638
rect 527 9582 613 9638
rect 669 9582 679 9638
rect 461 9496 679 9582
rect 461 9440 471 9496
rect 527 9440 613 9496
rect 669 9440 679 9496
rect 461 9354 679 9440
rect 461 9298 471 9354
rect 527 9298 613 9354
rect 669 9298 679 9354
rect 461 9212 679 9298
rect 461 9156 471 9212
rect 527 9156 613 9212
rect 669 9156 679 9212
rect 461 9070 679 9156
rect 461 9014 471 9070
rect 527 9014 613 9070
rect 669 9014 679 9070
rect 461 8928 679 9014
rect 461 8872 471 8928
rect 527 8872 613 8928
rect 669 8872 679 8928
rect 461 8786 679 8872
rect 461 8730 471 8786
rect 527 8730 613 8786
rect 669 8730 679 8786
rect 461 8644 679 8730
rect 461 8588 471 8644
rect 527 8588 613 8644
rect 669 8588 679 8644
rect 461 8502 679 8588
rect 461 8446 471 8502
rect 527 8446 613 8502
rect 669 8446 679 8502
rect 461 8360 679 8446
rect 461 8304 471 8360
rect 527 8304 613 8360
rect 669 8304 679 8360
rect 461 8218 679 8304
rect 461 8162 471 8218
rect 527 8162 613 8218
rect 669 8162 679 8218
rect 461 8076 679 8162
rect 461 8020 471 8076
rect 527 8020 613 8076
rect 669 8020 679 8076
rect 461 7934 679 8020
rect 461 7878 471 7934
rect 527 7878 613 7934
rect 669 7878 679 7934
rect 461 7792 679 7878
rect 461 7736 471 7792
rect 527 7736 613 7792
rect 669 7736 679 7792
rect 461 7650 679 7736
rect 461 7594 471 7650
rect 527 7594 613 7650
rect 669 7594 679 7650
rect 461 7508 679 7594
rect 461 7452 471 7508
rect 527 7452 613 7508
rect 669 7452 679 7508
rect 461 7366 679 7452
rect 461 7310 471 7366
rect 527 7310 613 7366
rect 669 7310 679 7366
rect 461 7224 679 7310
rect 461 7168 471 7224
rect 527 7168 613 7224
rect 669 7168 679 7224
rect 461 7082 679 7168
rect 461 7026 471 7082
rect 527 7026 613 7082
rect 669 7026 679 7082
rect 461 7016 679 7026
rect 11703 9922 11921 9932
rect 11703 9866 11713 9922
rect 11769 9866 11855 9922
rect 11911 9866 11921 9922
rect 11703 9780 11921 9866
rect 11703 9724 11713 9780
rect 11769 9724 11855 9780
rect 11911 9724 11921 9780
rect 11703 9638 11921 9724
rect 11703 9582 11713 9638
rect 11769 9582 11855 9638
rect 11911 9582 11921 9638
rect 11703 9496 11921 9582
rect 11703 9440 11713 9496
rect 11769 9440 11855 9496
rect 11911 9440 11921 9496
rect 11703 9354 11921 9440
rect 11703 9298 11713 9354
rect 11769 9298 11855 9354
rect 11911 9298 11921 9354
rect 11703 9212 11921 9298
rect 11703 9156 11713 9212
rect 11769 9156 11855 9212
rect 11911 9156 11921 9212
rect 11703 9070 11921 9156
rect 11703 9014 11713 9070
rect 11769 9014 11855 9070
rect 11911 9014 11921 9070
rect 11703 8928 11921 9014
rect 11703 8872 11713 8928
rect 11769 8872 11855 8928
rect 11911 8872 11921 8928
rect 11703 8786 11921 8872
rect 11703 8730 11713 8786
rect 11769 8730 11855 8786
rect 11911 8730 11921 8786
rect 11703 8644 11921 8730
rect 11703 8588 11713 8644
rect 11769 8588 11855 8644
rect 11911 8588 11921 8644
rect 11703 8502 11921 8588
rect 11703 8446 11713 8502
rect 11769 8446 11855 8502
rect 11911 8446 11921 8502
rect 11703 8360 11921 8446
rect 11703 8304 11713 8360
rect 11769 8304 11855 8360
rect 11911 8304 11921 8360
rect 11703 8218 11921 8304
rect 11703 8162 11713 8218
rect 11769 8162 11855 8218
rect 11911 8162 11921 8218
rect 11703 8076 11921 8162
rect 11703 8020 11713 8076
rect 11769 8020 11855 8076
rect 11911 8020 11921 8076
rect 11703 7934 11921 8020
rect 11703 7878 11713 7934
rect 11769 7878 11855 7934
rect 11911 7878 11921 7934
rect 11703 7792 11921 7878
rect 11703 7736 11713 7792
rect 11769 7736 11855 7792
rect 11911 7736 11921 7792
rect 11703 7650 11921 7736
rect 11703 7594 11713 7650
rect 11769 7594 11855 7650
rect 11911 7594 11921 7650
rect 11703 7508 11921 7594
rect 11703 7452 11713 7508
rect 11769 7452 11855 7508
rect 11911 7452 11921 7508
rect 11703 7366 11921 7452
rect 11703 7310 11713 7366
rect 11769 7310 11855 7366
rect 11911 7310 11921 7366
rect 11703 7224 11921 7310
rect 11703 7168 11713 7224
rect 11769 7168 11855 7224
rect 11911 7168 11921 7224
rect 11703 7082 11921 7168
rect 11703 7026 11713 7082
rect 11769 7026 11855 7082
rect 11911 7026 11921 7082
rect 11703 7016 11921 7026
rect 461 6740 679 6750
rect 461 6684 471 6740
rect 527 6684 613 6740
rect 669 6684 679 6740
rect 461 6598 679 6684
rect 461 6542 471 6598
rect 527 6542 613 6598
rect 669 6542 679 6598
rect 461 6456 679 6542
rect 461 6400 471 6456
rect 527 6400 613 6456
rect 669 6400 679 6456
rect 461 6314 679 6400
rect 461 6258 471 6314
rect 527 6258 613 6314
rect 669 6258 679 6314
rect 461 6172 679 6258
rect 461 6116 471 6172
rect 527 6116 613 6172
rect 669 6116 679 6172
rect 461 6030 679 6116
rect 461 5974 471 6030
rect 527 5974 613 6030
rect 669 5974 679 6030
rect 461 5888 679 5974
rect 461 5832 471 5888
rect 527 5832 613 5888
rect 669 5832 679 5888
rect 461 5746 679 5832
rect 461 5690 471 5746
rect 527 5690 613 5746
rect 669 5690 679 5746
rect 461 5604 679 5690
rect 461 5548 471 5604
rect 527 5548 613 5604
rect 669 5548 679 5604
rect 461 5462 679 5548
rect 461 5406 471 5462
rect 527 5406 613 5462
rect 669 5406 679 5462
rect 461 5320 679 5406
rect 461 5264 471 5320
rect 527 5264 613 5320
rect 669 5264 679 5320
rect 461 5178 679 5264
rect 461 5122 471 5178
rect 527 5122 613 5178
rect 669 5122 679 5178
rect 461 5036 679 5122
rect 461 4980 471 5036
rect 527 4980 613 5036
rect 669 4980 679 5036
rect 461 4894 679 4980
rect 461 4838 471 4894
rect 527 4838 613 4894
rect 669 4838 679 4894
rect 461 4752 679 4838
rect 461 4696 471 4752
rect 527 4696 613 4752
rect 669 4696 679 4752
rect 461 4610 679 4696
rect 461 4554 471 4610
rect 527 4554 613 4610
rect 669 4554 679 4610
rect 461 4468 679 4554
rect 461 4412 471 4468
rect 527 4412 613 4468
rect 669 4412 679 4468
rect 461 4326 679 4412
rect 461 4270 471 4326
rect 527 4270 613 4326
rect 669 4270 679 4326
rect 461 4184 679 4270
rect 461 4128 471 4184
rect 527 4128 613 4184
rect 669 4128 679 4184
rect 461 4042 679 4128
rect 461 3986 471 4042
rect 527 3986 613 4042
rect 669 3986 679 4042
rect 461 3900 679 3986
rect 461 3844 471 3900
rect 527 3844 613 3900
rect 669 3844 679 3900
rect 461 3834 679 3844
rect 11703 6740 11921 6750
rect 11703 6684 11713 6740
rect 11769 6684 11855 6740
rect 11911 6684 11921 6740
rect 11703 6598 11921 6684
rect 11703 6542 11713 6598
rect 11769 6542 11855 6598
rect 11911 6542 11921 6598
rect 11703 6456 11921 6542
rect 11703 6400 11713 6456
rect 11769 6400 11855 6456
rect 11911 6400 11921 6456
rect 11703 6314 11921 6400
rect 11703 6258 11713 6314
rect 11769 6258 11855 6314
rect 11911 6258 11921 6314
rect 11703 6172 11921 6258
rect 11703 6116 11713 6172
rect 11769 6116 11855 6172
rect 11911 6116 11921 6172
rect 11703 6030 11921 6116
rect 11703 5974 11713 6030
rect 11769 5974 11855 6030
rect 11911 5974 11921 6030
rect 11703 5888 11921 5974
rect 11703 5832 11713 5888
rect 11769 5832 11855 5888
rect 11911 5832 11921 5888
rect 11703 5746 11921 5832
rect 11703 5690 11713 5746
rect 11769 5690 11855 5746
rect 11911 5690 11921 5746
rect 11703 5604 11921 5690
rect 11703 5548 11713 5604
rect 11769 5548 11855 5604
rect 11911 5548 11921 5604
rect 11703 5462 11921 5548
rect 11703 5406 11713 5462
rect 11769 5406 11855 5462
rect 11911 5406 11921 5462
rect 11703 5320 11921 5406
rect 11703 5264 11713 5320
rect 11769 5264 11855 5320
rect 11911 5264 11921 5320
rect 11703 5178 11921 5264
rect 11703 5122 11713 5178
rect 11769 5122 11855 5178
rect 11911 5122 11921 5178
rect 11703 5036 11921 5122
rect 11703 4980 11713 5036
rect 11769 4980 11855 5036
rect 11911 4980 11921 5036
rect 11703 4894 11921 4980
rect 11703 4838 11713 4894
rect 11769 4838 11855 4894
rect 11911 4838 11921 4894
rect 11703 4752 11921 4838
rect 11703 4696 11713 4752
rect 11769 4696 11855 4752
rect 11911 4696 11921 4752
rect 11703 4610 11921 4696
rect 11703 4554 11713 4610
rect 11769 4554 11855 4610
rect 11911 4554 11921 4610
rect 11703 4468 11921 4554
rect 11703 4412 11713 4468
rect 11769 4412 11855 4468
rect 11911 4412 11921 4468
rect 11703 4326 11921 4412
rect 11703 4270 11713 4326
rect 11769 4270 11855 4326
rect 11911 4270 11921 4326
rect 11703 4184 11921 4270
rect 11703 4128 11713 4184
rect 11769 4128 11855 4184
rect 11911 4128 11921 4184
rect 11703 4042 11921 4128
rect 11703 3986 11713 4042
rect 11769 3986 11855 4042
rect 11911 3986 11921 4042
rect 11703 3900 11921 3986
rect 11703 3844 11713 3900
rect 11769 3844 11855 3900
rect 11911 3844 11921 3900
rect 11703 3834 11921 3844
rect 461 3522 679 3532
rect 461 3466 471 3522
rect 527 3466 613 3522
rect 669 3466 679 3522
rect 461 3380 679 3466
rect 461 3324 471 3380
rect 527 3324 613 3380
rect 669 3324 679 3380
rect 461 3238 679 3324
rect 461 3182 471 3238
rect 527 3182 613 3238
rect 669 3182 679 3238
rect 461 3096 679 3182
rect 461 3040 471 3096
rect 527 3040 613 3096
rect 669 3040 679 3096
rect 461 3030 679 3040
rect 11703 3522 11921 3532
rect 11703 3466 11713 3522
rect 11769 3466 11855 3522
rect 11911 3466 11921 3522
rect 11703 3380 11921 3466
rect 11703 3324 11713 3380
rect 11769 3324 11855 3380
rect 11911 3324 11921 3380
rect 11703 3238 11921 3324
rect 11703 3182 11713 3238
rect 11769 3182 11855 3238
rect 11911 3182 11921 3238
rect 11703 3096 11921 3182
rect 11703 3040 11713 3096
rect 11769 3040 11855 3096
rect 11911 3040 11921 3096
rect 11703 3030 11921 3040
rect 442 2317 802 2327
rect 442 2261 452 2317
rect 508 2261 594 2317
rect 650 2261 736 2317
rect 792 2261 802 2317
rect 442 2175 802 2261
rect 442 2119 452 2175
rect 508 2119 594 2175
rect 650 2119 736 2175
rect 792 2119 802 2175
rect 442 2033 802 2119
rect 442 1977 452 2033
rect 508 1977 594 2033
rect 650 1977 736 2033
rect 792 1977 802 2033
rect 442 1891 802 1977
rect 442 1835 452 1891
rect 508 1835 594 1891
rect 650 1835 736 1891
rect 792 1835 802 1891
rect 442 1749 802 1835
rect 442 1693 452 1749
rect 508 1693 594 1749
rect 650 1693 736 1749
rect 792 1693 802 1749
rect 442 1607 802 1693
rect 442 1551 452 1607
rect 508 1551 594 1607
rect 650 1551 736 1607
rect 792 1551 802 1607
rect 442 1465 802 1551
rect 442 1409 452 1465
rect 508 1409 594 1465
rect 650 1409 736 1465
rect 792 1409 802 1465
rect 442 1323 802 1409
rect 442 1267 452 1323
rect 508 1267 594 1323
rect 650 1267 736 1323
rect 792 1267 802 1323
rect 442 1181 802 1267
rect 442 1125 452 1181
rect 508 1125 594 1181
rect 650 1125 736 1181
rect 792 1125 802 1181
rect 442 1039 802 1125
rect 442 983 452 1039
rect 508 983 594 1039
rect 650 983 736 1039
rect 792 983 802 1039
rect 442 897 802 983
rect 442 841 452 897
rect 508 841 594 897
rect 650 841 736 897
rect 792 841 802 897
rect 442 755 802 841
rect 442 699 452 755
rect 508 699 594 755
rect 650 699 736 755
rect 792 699 802 755
rect 442 689 802 699
rect 11571 2317 11931 2327
rect 11571 2261 11581 2317
rect 11637 2261 11723 2317
rect 11779 2261 11865 2317
rect 11921 2261 11931 2317
rect 11571 2175 11931 2261
rect 11571 2119 11581 2175
rect 11637 2119 11723 2175
rect 11779 2119 11865 2175
rect 11921 2119 11931 2175
rect 11571 2033 11931 2119
rect 11571 1977 11581 2033
rect 11637 1977 11723 2033
rect 11779 1977 11865 2033
rect 11921 1977 11931 2033
rect 11571 1891 11931 1977
rect 11571 1835 11581 1891
rect 11637 1835 11723 1891
rect 11779 1835 11865 1891
rect 11921 1835 11931 1891
rect 11571 1749 11931 1835
rect 11571 1693 11581 1749
rect 11637 1693 11723 1749
rect 11779 1693 11865 1749
rect 11921 1693 11931 1749
rect 11571 1607 11931 1693
rect 11571 1551 11581 1607
rect 11637 1551 11723 1607
rect 11779 1551 11865 1607
rect 11921 1551 11931 1607
rect 11571 1465 11931 1551
rect 11571 1409 11581 1465
rect 11637 1409 11723 1465
rect 11779 1409 11865 1465
rect 11921 1409 11931 1465
rect 11571 1323 11931 1409
rect 11571 1267 11581 1323
rect 11637 1267 11723 1323
rect 11779 1267 11865 1323
rect 11921 1267 11931 1323
rect 11571 1181 11931 1267
rect 11571 1125 11581 1181
rect 11637 1125 11723 1181
rect 11779 1125 11865 1181
rect 11921 1125 11931 1181
rect 11571 1039 11931 1125
rect 11571 983 11581 1039
rect 11637 983 11723 1039
rect 11779 983 11865 1039
rect 11921 983 11931 1039
rect 11571 897 11931 983
rect 11571 841 11581 897
rect 11637 841 11723 897
rect 11779 841 11865 897
rect 11921 841 11931 897
rect 11571 755 11931 841
rect 11571 699 11581 755
rect 11637 699 11723 755
rect 11779 699 11865 755
rect 11921 699 11931 755
rect 11571 689 11931 699
rect 12860 356 13078 366
rect 12860 300 12870 356
rect 12926 300 13012 356
rect 13068 300 13078 356
rect -727 288 -509 298
rect -727 232 -717 288
rect -661 232 -575 288
rect -519 232 -509 288
rect -727 146 -509 232
rect -727 90 -717 146
rect -661 90 -575 146
rect -519 90 -509 146
rect -727 4 -509 90
rect -727 -52 -717 4
rect -661 -52 -575 4
rect -519 -52 -509 4
rect -727 -138 -509 -52
rect -727 -194 -717 -138
rect -661 -194 -575 -138
rect -519 -194 -509 -138
rect -727 -280 -509 -194
rect -727 -336 -717 -280
rect -661 -336 -575 -280
rect -519 -336 -509 -280
rect -727 -422 -509 -336
rect -727 -478 -717 -422
rect -661 -478 -575 -422
rect -519 -478 -509 -422
rect -727 -564 -509 -478
rect -727 -620 -717 -564
rect -661 -620 -575 -564
rect -519 -620 -509 -564
rect -727 -706 -509 -620
rect -727 -762 -717 -706
rect -661 -762 -575 -706
rect -519 -762 -509 -706
rect -727 -848 -509 -762
rect -727 -904 -717 -848
rect -661 -904 -575 -848
rect -519 -904 -509 -848
rect -727 -914 -509 -904
rect 12860 214 13078 300
rect 12860 158 12870 214
rect 12926 158 13012 214
rect 13068 158 13078 214
rect 12860 72 13078 158
rect 12860 16 12870 72
rect 12926 16 13012 72
rect 13068 16 13078 72
rect 12860 -70 13078 16
rect 12860 -126 12870 -70
rect 12926 -126 13012 -70
rect 13068 -126 13078 -70
rect 12860 -212 13078 -126
rect 12860 -268 12870 -212
rect 12926 -268 13012 -212
rect 13068 -268 13078 -212
rect 12860 -354 13078 -268
rect 12860 -410 12870 -354
rect 12926 -410 13012 -354
rect 13068 -410 13078 -354
rect 12860 -496 13078 -410
rect 12860 -552 12870 -496
rect 12926 -552 13012 -496
rect 13068 -552 13078 -496
rect 12860 -638 13078 -552
rect 12860 -694 12870 -638
rect 12926 -694 13012 -638
rect 13068 -694 13078 -638
rect 12860 -780 13078 -694
rect 12860 -836 12870 -780
rect 12926 -836 13012 -780
rect 13068 -836 13078 -780
rect 12860 -922 13078 -836
rect 12860 -978 12870 -922
rect 12926 -978 13012 -922
rect 13068 -978 13078 -922
rect 12860 -988 13078 -978
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_0
timestamp 1764353313
transform -1 0 6347 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_1
timestamp 1764353313
transform -1 0 11651 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_2
timestamp 1764353313
transform 1 0 6035 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_3
timestamp 1764353313
transform 1 0 731 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_0
timestamp 1764353313
transform -1 0 4579 0 1 2840
box 0 12 1196 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_1
timestamp 1764353313
transform -1 0 9883 0 1 2840
box 0 12 1196 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_2
timestamp 1764353313
transform 1 0 2499 0 1 2840
box 0 12 1196 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_3
timestamp 1764353313
transform 1 0 7803 0 1 2840
box 0 12 1196 8252
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_0
timestamp 1764353313
transform -1 0 11573 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_1
timestamp 1764353313
transform 1 0 2577 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_2
timestamp 1764353313
transform 1 0 4345 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_3
timestamp 1764353313
transform 1 0 6113 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_4
timestamp 1764353313
transform 1 0 7881 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_5
timestamp 1764353313
transform 1 0 9649 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_6
timestamp 1764353313
transform 1 0 809 0 1 2972
box -44 0 1584 8000
<< properties >>
string GDS_END 13422302
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 12687920
<< end >>
