magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< obsm1 >>
rect -32 13108 1032 69957
<< obsm2 >>
rect 0 13622 1000 69616
<< obsm3 >>
rect 0 49200 1000 65000
<< obsm4 >>
rect 0 49200 1000 65000
<< metal5 >>
rect 0 63600 1000 65000
rect 0 49200 1000 50600
<< labels >>
rlabel metal5 s 0 63600 1000 65000 6 VSS
port 1 nsew ground bidirectional
rlabel metal5 s 0 49200 1000 50600 6 VSS
port 1 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 14144420
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 14136094
<< end >>
