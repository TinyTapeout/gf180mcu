magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< psubdiff >>
rect 13097 70975 69968 71000
rect 13097 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69968 70975
rect 13097 70871 69968 70929
rect 13097 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69968 70871
rect 13097 70803 69968 70825
rect 13097 70767 13291 70803
rect 13097 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13291 70767
rect 13097 70663 13291 70721
rect 13097 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13291 70663
rect 13097 70559 13291 70617
rect 13097 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13291 70559
rect 13097 70455 13291 70513
rect 13097 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13291 70455
rect 13097 70351 13291 70409
rect 13097 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13291 70351
rect 13097 70247 13291 70305
rect 13097 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13291 70247
rect 13097 70143 13291 70201
rect 13097 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13291 70143
rect 13097 70039 13291 70097
rect 13097 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13291 70039
rect 13097 69935 13291 69993
rect 13097 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13291 69935
rect 13097 69831 13291 69889
rect 13097 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13291 69831
rect 13097 69727 13291 69785
rect 69774 70720 69968 70803
rect 69774 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69968 70720
rect 69774 70616 69968 70674
rect 69774 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69968 70616
rect 69774 70512 69968 70570
rect 69774 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69968 70512
rect 69774 70408 69968 70466
rect 69774 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69968 70408
rect 69774 70304 69968 70362
rect 69774 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69968 70304
rect 69774 70200 69968 70258
rect 69774 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69968 70200
rect 69774 70096 69968 70154
rect 69774 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69968 70096
rect 69774 69968 69968 70050
rect 69774 69946 71000 69968
rect 69774 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69774 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69774 69842 71000 69862
rect 69774 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69774 69774 70824 69796
rect 13097 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13291 69727
rect 13097 69623 13291 69681
rect 13097 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13291 69623
rect 13097 69519 13291 69577
rect 13097 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13291 69519
rect 13097 69415 13291 69473
rect 13097 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13291 69415
rect 13097 69311 13291 69369
rect 13097 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13291 69311
rect 13097 69207 13291 69265
rect 13097 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13291 69207
rect 13097 69103 13291 69161
rect 13097 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13291 69103
rect 13097 68999 13291 69057
rect 13097 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13291 68999
rect 13097 68895 13291 68953
rect 13097 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13291 68895
rect 13097 68791 13291 68849
rect 13097 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13291 68791
rect 13097 68687 13291 68745
rect 13097 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13291 68687
rect 13097 68583 13291 68641
rect 13097 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13291 68583
rect 13097 68479 13291 68537
rect 13097 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13291 68479
rect 13097 68375 13291 68433
rect 13097 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13291 68375
rect 13097 68271 13291 68329
rect 13097 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13291 68271
rect 13097 68167 13291 68225
rect 13097 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13291 68167
rect 13097 68063 13291 68121
rect 13097 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13291 68063
rect 13097 67959 13291 68017
rect 13097 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13291 67959
rect 13097 67855 13291 67913
rect 13097 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13291 67855
rect 13097 67751 13291 67809
rect 13097 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13291 67751
rect 13097 67647 13291 67705
rect 13097 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13291 67647
rect 13097 67543 13291 67601
rect 13097 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13291 67543
rect 13097 67439 13291 67497
rect 13097 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13291 67439
rect 13097 67335 13291 67393
rect 13097 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13291 67335
rect 13097 67231 13291 67289
rect 13097 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13291 67231
rect 13097 67127 13291 67185
rect 13097 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13291 67127
rect 13097 67023 13291 67081
rect 13097 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13291 67023
rect 13097 66919 13291 66977
rect 13097 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13291 66919
rect 13097 66815 13291 66873
rect 13097 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13291 66815
rect 13097 66711 13291 66769
rect 13097 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13291 66711
rect 13097 66607 13291 66665
rect 13097 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13291 66607
rect 13097 66503 13291 66561
rect 13097 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13291 66503
rect 13097 66399 13291 66457
rect 13097 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13291 66399
rect 13097 66295 13291 66353
rect 13097 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13291 66295
rect 13097 66191 13291 66249
rect 13097 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13291 66191
rect 13097 66087 13291 66145
rect 13097 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13291 66087
rect 13097 65983 13291 66041
rect 13097 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13291 65983
rect 13097 65879 13291 65937
rect 13097 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13291 65879
rect 13097 65775 13291 65833
rect 13097 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13291 65775
rect 13097 65671 13291 65729
rect 13097 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13291 65671
rect 13097 65567 13291 65625
rect 13097 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13291 65567
rect 13097 65463 13291 65521
rect 13097 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13291 65463
rect 13097 65359 13291 65417
rect 13097 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13291 65359
rect 13097 65255 13291 65313
rect 13097 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13291 65255
rect 13097 65151 13291 65209
rect 13097 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13291 65151
rect 13097 65047 13291 65105
rect 13097 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13291 65047
rect 13097 64943 13291 65001
rect 13097 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13291 64943
rect 13097 64839 13291 64897
rect 13097 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13291 64839
rect 13097 64735 13291 64793
rect 13097 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13291 64735
rect 13097 64631 13291 64689
rect 13097 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13291 64631
rect 13097 64527 13291 64585
rect 13097 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13291 64527
rect 13097 64423 13291 64481
rect 13097 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13291 64423
rect 13097 64319 13291 64377
rect 13097 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13291 64319
rect 13097 64215 13291 64273
rect 13097 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13291 64215
rect 13097 64111 13291 64169
rect 13097 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13291 64111
rect 13097 64007 13291 64065
rect 13097 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13291 64007
rect 13097 63903 13291 63961
rect 13097 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13291 63903
rect 13097 63799 13291 63857
rect 13097 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13291 63799
rect 13097 63695 13291 63753
rect 13097 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13291 63695
rect 13097 63591 13291 63649
rect 13097 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13291 63591
rect 13097 63487 13291 63545
rect 13097 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13291 63487
rect 13097 63383 13291 63441
rect 13097 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13291 63383
rect 13097 63279 13291 63337
rect 13097 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13291 63279
rect 13097 63175 13291 63233
rect 13097 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13291 63175
rect 13097 63071 13291 63129
rect 13097 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13291 63071
rect 13097 62967 13291 63025
rect 13097 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13291 62967
rect 13097 62863 13291 62921
rect 13097 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13291 62863
rect 13097 62759 13291 62817
rect 13097 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13291 62759
rect 13097 62655 13291 62713
rect 13097 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13291 62655
rect 13097 62551 13291 62609
rect 13097 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13291 62551
rect 13097 62447 13291 62505
rect 13097 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13291 62447
rect 13097 62343 13291 62401
rect 13097 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13291 62343
rect 13097 62239 13291 62297
rect 13097 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13291 62239
rect 13097 62135 13291 62193
rect 13097 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13291 62135
rect 13097 62031 13291 62089
rect 13097 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13291 62031
rect 13097 61927 13291 61985
rect 13097 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13291 61927
rect 13097 61823 13291 61881
rect 13097 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13291 61823
rect 13097 61719 13291 61777
rect 13097 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13291 61719
rect 13097 61615 13291 61673
rect 13097 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13291 61615
rect 13097 61511 13291 61569
rect 13097 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13291 61511
rect 13097 61407 13291 61465
rect 13097 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13291 61407
rect 13097 61303 13291 61361
rect 13097 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13291 61303
rect 13097 61199 13291 61257
rect 13097 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13291 61199
rect 13097 61095 13291 61153
rect 13097 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13291 61095
rect 13097 60991 13291 61049
rect 13097 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13291 60991
rect 13097 60887 13291 60945
rect 13097 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13291 60887
rect 13097 60783 13291 60841
rect 13097 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13291 60783
rect 13097 60679 13291 60737
rect 13097 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13291 60679
rect 13097 60575 13291 60633
rect 13097 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13291 60575
rect 13097 60471 13291 60529
rect 13097 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13291 60471
rect 13097 60367 13291 60425
rect 13097 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13291 60367
rect 13097 60263 13291 60321
rect 13097 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13291 60263
rect 13097 60159 13291 60217
rect 13097 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13291 60159
rect 13097 60055 13291 60113
rect 13097 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13291 60055
rect 13097 59951 13291 60009
rect 13097 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13291 59951
rect 13097 59847 13291 59905
rect 13097 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13291 59847
rect 13097 59743 13291 59801
rect 13097 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13291 59743
rect 13097 59639 13291 59697
rect 13097 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13291 59639
rect 13097 59535 13291 59593
rect 13097 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13291 59535
rect 13097 59431 13291 59489
rect 13097 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13291 59431
rect 13097 59327 13291 59385
rect 13097 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13291 59327
rect 13097 59223 13291 59281
rect 13097 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13291 59223
rect 13097 59119 13291 59177
rect 13097 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13291 59119
rect 13097 59015 13291 59073
rect 13097 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13291 59015
rect 13097 58911 13291 58969
rect 13097 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13291 58911
rect 13097 58807 13291 58865
rect 13097 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13291 58807
rect 13097 58703 13291 58761
rect 13097 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13291 58703
rect 13097 58599 13291 58657
rect 13097 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13291 58599
rect 13097 58495 13291 58553
rect 13097 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13291 58495
rect 13097 58391 13291 58449
rect 13097 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13291 58391
rect 13097 58287 13291 58345
rect 13097 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13291 58287
rect 13097 58183 13291 58241
rect 13097 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13291 58183
rect 13097 58079 13291 58137
rect 13097 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13291 58079
rect 13097 57975 13291 58033
rect 13097 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13291 57975
rect 13097 57871 13291 57929
rect 13097 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13291 57871
rect 13097 57767 13291 57825
rect 13097 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13291 57767
rect 13097 57663 13291 57721
rect 13097 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13291 57663
rect 13097 57559 13291 57617
rect 13097 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13291 57559
rect 13097 57455 13291 57513
rect 13097 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13291 57455
rect 13097 57351 13291 57409
rect 13097 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13291 57351
rect 13097 57247 13291 57305
rect 13097 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13291 57247
rect 13097 57143 13291 57201
rect 13097 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13291 57143
rect 13097 57039 13291 57097
rect 13097 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13291 57039
rect 13097 56935 13291 56993
rect 13097 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13291 56935
rect 13097 56831 13291 56889
rect 13097 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13291 56831
rect 13097 56727 13291 56785
rect 13097 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13291 56727
rect 13097 56623 13291 56681
rect 13097 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13291 56623
rect 13097 56519 13291 56577
rect 13097 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13291 56519
rect 13097 56415 13291 56473
rect 13097 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13291 56415
rect 13097 56311 13291 56369
rect 13097 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13291 56311
rect 13097 56207 13291 56265
rect 13097 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13291 56207
rect 13097 56103 13291 56161
rect 13097 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13291 56103
rect 13097 55999 13291 56057
rect 13097 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13291 55999
rect 13097 55895 13291 55953
rect 13097 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13291 55895
rect 13097 55791 13291 55849
rect 13097 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13291 55791
rect 13097 55687 13291 55745
rect 13097 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13291 55687
rect 13097 55583 13291 55641
rect 13097 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13291 55583
rect 13097 55479 13291 55537
rect 13097 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13291 55479
rect 13097 55375 13291 55433
rect 13097 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13291 55375
rect 13097 55271 13291 55329
rect 13097 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13291 55271
rect 13097 55167 13291 55225
rect 13097 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13291 55167
rect 13097 55063 13291 55121
rect 13097 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13291 55063
rect 13097 54959 13291 55017
rect 13097 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13291 54959
rect 13097 54855 13291 54913
rect 13097 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13291 54855
rect 13097 54751 13291 54809
rect 13097 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13291 54751
rect 13097 54647 13291 54705
rect 13097 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13291 54647
rect 13097 54543 13291 54601
rect 13097 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13291 54543
rect 13097 54439 13291 54497
rect 13097 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13291 54439
rect 13097 54335 13291 54393
rect 13097 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13291 54335
rect 13097 54231 13291 54289
rect 13097 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13291 54231
rect 13097 54127 13291 54185
rect 13097 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13291 54127
rect 13097 54023 13291 54081
rect 13097 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13291 54023
rect 13097 53919 13291 53977
rect 13097 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13291 53919
rect 13097 53815 13291 53873
rect 13097 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13291 53815
rect 13097 53711 13291 53769
rect 13097 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13291 53711
rect 13097 53607 13291 53665
rect 13097 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13291 53607
rect 13097 53503 13291 53561
rect 13097 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13291 53503
rect 13097 53399 13291 53457
rect 13097 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13291 53399
rect 13097 53295 13291 53353
rect 13097 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13291 53295
rect 13097 53191 13291 53249
rect 13097 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13291 53191
rect 13097 53087 13291 53145
rect 13097 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13291 53087
rect 13097 52983 13291 53041
rect 13097 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13291 52983
rect 13097 52879 13291 52937
rect 13097 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13291 52879
rect 13097 52775 13291 52833
rect 13097 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13291 52775
rect 13097 52671 13291 52729
rect 13097 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13291 52671
rect 13097 52567 13291 52625
rect 13097 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13291 52567
rect 13097 52463 13291 52521
rect 13097 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13291 52463
rect 13097 52359 13291 52417
rect 13097 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13291 52359
rect 13097 52255 13291 52313
rect 13097 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13291 52255
rect 13097 52151 13291 52209
rect 13097 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13291 52151
rect 13097 52047 13291 52105
rect 13097 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13291 52047
rect 13097 51943 13291 52001
rect 13097 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13291 51943
rect 13097 51839 13291 51897
rect 13097 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13291 51839
rect 13097 51735 13291 51793
rect 13097 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13291 51735
rect 13097 51631 13291 51689
rect 13097 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13291 51631
rect 13097 51527 13291 51585
rect 13097 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13291 51527
rect 13097 51423 13291 51481
rect 13097 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13291 51423
rect 13097 51319 13291 51377
rect 13097 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13291 51319
rect 13097 51215 13291 51273
rect 13097 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13291 51215
rect 13097 51111 13291 51169
rect 13097 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13291 51111
rect 13097 51007 13291 51065
rect 13097 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13291 51007
rect 13097 50903 13291 50961
rect 13097 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13291 50903
rect 13097 50799 13291 50857
rect 13097 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13291 50799
rect 13097 50695 13291 50753
rect 13097 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13291 50695
rect 13097 50591 13291 50649
rect 13097 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13291 50591
rect 13097 50487 13291 50545
rect 13097 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13291 50487
rect 13097 50383 13291 50441
rect 13097 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13291 50383
rect 13097 50279 13291 50337
rect 13097 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13291 50279
rect 13097 50175 13291 50233
rect 13097 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13291 50175
rect 13097 50071 13291 50129
rect 13097 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13291 50071
rect 13097 49967 13291 50025
rect 13097 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13291 49967
rect 13097 49863 13291 49921
rect 13097 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13291 49863
rect 13097 49759 13291 49817
rect 13097 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13291 49759
rect 13097 49655 13291 49713
rect 13097 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13291 49655
rect 13097 49551 13291 49609
rect 13097 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13291 49551
rect 13097 49447 13291 49505
rect 13097 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13291 49447
rect 13097 49343 13291 49401
rect 13097 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13291 49343
rect 13097 49239 13291 49297
rect 13097 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13291 49239
rect 13097 49135 13291 49193
rect 13097 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13291 49135
rect 13097 49031 13291 49089
rect 13097 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13291 49031
rect 13097 48927 13291 48985
rect 13097 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13291 48927
rect 13097 48823 13291 48881
rect 13097 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13291 48823
rect 13097 48719 13291 48777
rect 13097 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13291 48719
rect 13097 48615 13291 48673
rect 13097 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13291 48615
rect 13097 48511 13291 48569
rect 13097 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13291 48511
rect 13097 48407 13291 48465
rect 13097 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13291 48407
rect 13097 48303 13291 48361
rect 13097 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13291 48303
rect 13097 48199 13291 48257
rect 13097 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13291 48199
rect 13097 48095 13291 48153
rect 13097 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13291 48095
rect 13097 47991 13291 48049
rect 13097 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13291 47991
rect 13097 47887 13291 47945
rect 13097 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13291 47887
rect 13097 47783 13291 47841
rect 13097 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13291 47783
rect 13097 47679 13291 47737
rect 13097 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13291 47679
rect 13097 47575 13291 47633
rect 13097 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13291 47575
rect 13097 47471 13291 47529
rect 13097 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13291 47471
rect 13097 47367 13291 47425
rect 13097 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13291 47367
rect 13097 47263 13291 47321
rect 13097 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13291 47263
rect 13097 47159 13291 47217
rect 13097 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13291 47159
rect 13097 47055 13291 47113
rect 13097 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13291 47055
rect 13097 46951 13291 47009
rect 13097 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13291 46951
rect 13097 46847 13291 46905
rect 13097 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13291 46847
rect 13097 46743 13291 46801
rect 13097 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13291 46743
rect 13097 46639 13291 46697
rect 13097 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13291 46639
rect 13097 46535 13291 46593
rect 13097 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13291 46535
rect 13097 46431 13291 46489
rect 13097 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13291 46431
rect 13097 46327 13291 46385
rect 13097 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13291 46327
rect 13097 46223 13291 46281
rect 13097 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13291 46223
rect 13097 46119 13291 46177
rect 13097 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13291 46119
rect 13097 46015 13291 46073
rect 13097 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13291 46015
rect 13097 45911 13291 45969
rect 13097 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13291 45911
rect 13097 45807 13291 45865
rect 13097 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13291 45807
rect 13097 45703 13291 45761
rect 13097 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13291 45703
rect 13097 45599 13291 45657
rect 13097 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13291 45599
rect 13097 45495 13291 45553
rect 13097 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13291 45495
rect 13097 45391 13291 45449
rect 13097 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13291 45391
rect 13097 45287 13291 45345
rect 13097 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13291 45287
rect 13097 45183 13291 45241
rect 13097 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13291 45183
rect 13097 45079 13291 45137
rect 13097 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13291 45079
rect 13097 44921 13291 45033
rect 70802 69758 70824 69774
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70802 69700 71000 69758
rect 70802 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70802 69596 71000 69654
rect 70802 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70802 69492 71000 69550
rect 70802 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70802 69388 71000 69446
rect 70802 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70802 69284 71000 69342
rect 70802 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70802 69180 71000 69238
rect 70802 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70802 69076 71000 69134
rect 70802 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70802 68972 71000 69030
rect 70802 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70802 68868 71000 68926
rect 70802 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70802 68764 71000 68822
rect 70802 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70802 68660 71000 68718
rect 70802 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70802 68556 71000 68614
rect 70802 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70802 68452 71000 68510
rect 70802 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70802 68348 71000 68406
rect 70802 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70802 68244 71000 68302
rect 70802 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70802 68140 71000 68198
rect 70802 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70802 68036 71000 68094
rect 70802 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70802 67932 71000 67990
rect 70802 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70802 67828 71000 67886
rect 70802 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70802 67724 71000 67782
rect 70802 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70802 67620 71000 67678
rect 70802 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70802 67516 71000 67574
rect 70802 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70802 67412 71000 67470
rect 70802 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70802 67308 71000 67366
rect 70802 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70802 67204 71000 67262
rect 70802 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70802 67100 71000 67158
rect 70802 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70802 66996 71000 67054
rect 70802 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70802 66892 71000 66950
rect 70802 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70802 66788 71000 66846
rect 70802 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70802 66684 71000 66742
rect 70802 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70802 66580 71000 66638
rect 70802 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70802 66476 71000 66534
rect 70802 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70802 66372 71000 66430
rect 70802 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70802 66268 71000 66326
rect 70802 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70802 66164 71000 66222
rect 70802 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70802 66060 71000 66118
rect 70802 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70802 65956 71000 66014
rect 70802 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70802 65852 71000 65910
rect 70802 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70802 65748 71000 65806
rect 70802 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70802 65644 71000 65702
rect 70802 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70802 65540 71000 65598
rect 70802 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70802 65436 71000 65494
rect 70802 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70802 65332 71000 65390
rect 70802 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70802 65228 71000 65286
rect 70802 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70802 65124 71000 65182
rect 70802 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70802 65020 71000 65078
rect 70802 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70802 64916 71000 64974
rect 70802 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70802 64812 71000 64870
rect 70802 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70802 64708 71000 64766
rect 70802 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70802 64604 71000 64662
rect 70802 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70802 64500 71000 64558
rect 70802 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70802 64396 71000 64454
rect 70802 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70802 64292 71000 64350
rect 70802 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70802 64188 71000 64246
rect 70802 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70802 64084 71000 64142
rect 70802 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70802 63980 71000 64038
rect 70802 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70802 63876 71000 63934
rect 70802 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70802 63772 71000 63830
rect 70802 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70802 63668 71000 63726
rect 70802 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70802 63564 71000 63622
rect 70802 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70802 63460 71000 63518
rect 70802 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70802 63356 71000 63414
rect 70802 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70802 63252 71000 63310
rect 70802 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70802 63148 71000 63206
rect 70802 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70802 63044 71000 63102
rect 70802 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70802 62940 71000 62998
rect 70802 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70802 62836 71000 62894
rect 70802 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70802 62732 71000 62790
rect 70802 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70802 62628 71000 62686
rect 70802 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70802 62524 71000 62582
rect 70802 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70802 62420 71000 62478
rect 70802 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70802 62316 71000 62374
rect 70802 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70802 62212 71000 62270
rect 70802 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70802 62108 71000 62166
rect 70802 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70802 62004 71000 62062
rect 70802 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70802 61900 71000 61958
rect 70802 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70802 61796 71000 61854
rect 70802 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70802 61692 71000 61750
rect 70802 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70802 61588 71000 61646
rect 70802 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70802 61484 71000 61542
rect 70802 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70802 61380 71000 61438
rect 70802 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70802 61276 71000 61334
rect 70802 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70802 61172 71000 61230
rect 70802 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70802 61068 71000 61126
rect 70802 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70802 60964 71000 61022
rect 70802 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70802 60860 71000 60918
rect 70802 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70802 60756 71000 60814
rect 70802 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70802 60652 71000 60710
rect 70802 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70802 60548 71000 60606
rect 70802 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70802 60444 71000 60502
rect 70802 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70802 60340 71000 60398
rect 70802 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70802 60236 71000 60294
rect 70802 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70802 60132 71000 60190
rect 70802 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70802 60028 71000 60086
rect 70802 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70802 59924 71000 59982
rect 70802 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70802 59820 71000 59878
rect 70802 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70802 59716 71000 59774
rect 70802 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70802 59612 71000 59670
rect 70802 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70802 59508 71000 59566
rect 70802 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70802 59404 71000 59462
rect 70802 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70802 59300 71000 59358
rect 70802 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70802 59196 71000 59254
rect 70802 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70802 59092 71000 59150
rect 70802 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70802 58988 71000 59046
rect 70802 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70802 58884 71000 58942
rect 70802 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70802 58780 71000 58838
rect 70802 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70802 58676 71000 58734
rect 70802 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70802 58572 71000 58630
rect 70802 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70802 58468 71000 58526
rect 70802 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70802 58364 71000 58422
rect 70802 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70802 58260 71000 58318
rect 70802 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70802 58156 71000 58214
rect 70802 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70802 58052 71000 58110
rect 70802 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70802 57948 71000 58006
rect 70802 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70802 57844 71000 57902
rect 70802 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70802 57740 71000 57798
rect 70802 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70802 57636 71000 57694
rect 70802 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70802 57532 71000 57590
rect 70802 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70802 57428 71000 57486
rect 70802 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70802 57324 71000 57382
rect 70802 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70802 57220 71000 57278
rect 70802 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70802 57116 71000 57174
rect 70802 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70802 57012 71000 57070
rect 70802 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70802 56908 71000 56966
rect 70802 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70802 56804 71000 56862
rect 70802 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70802 56700 71000 56758
rect 70802 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70802 56596 71000 56654
rect 70802 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70802 56492 71000 56550
rect 70802 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70802 56388 71000 56446
rect 70802 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70802 56284 71000 56342
rect 70802 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70802 56180 71000 56238
rect 70802 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70802 56076 71000 56134
rect 70802 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70802 55972 71000 56030
rect 70802 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70802 55868 71000 55926
rect 70802 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70802 55764 71000 55822
rect 70802 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70802 55660 71000 55718
rect 70802 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70802 55556 71000 55614
rect 70802 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70802 55452 71000 55510
rect 70802 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70802 55348 71000 55406
rect 70802 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70802 55244 71000 55302
rect 70802 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70802 55140 71000 55198
rect 70802 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70802 55036 71000 55094
rect 70802 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70802 54932 71000 54990
rect 70802 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70802 54828 71000 54886
rect 70802 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70802 54724 71000 54782
rect 70802 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70802 54620 71000 54678
rect 70802 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70802 54516 71000 54574
rect 70802 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70802 54412 71000 54470
rect 70802 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70802 54308 71000 54366
rect 70802 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70802 54204 71000 54262
rect 70802 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70802 54100 71000 54158
rect 70802 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70802 53996 71000 54054
rect 70802 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70802 53892 71000 53950
rect 70802 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70802 53788 71000 53846
rect 70802 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70802 53684 71000 53742
rect 70802 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70802 53580 71000 53638
rect 70802 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70802 53476 71000 53534
rect 70802 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70802 53372 71000 53430
rect 70802 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70802 53268 71000 53326
rect 70802 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70802 53164 71000 53222
rect 70802 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70802 53060 71000 53118
rect 70802 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70802 52956 71000 53014
rect 70802 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70802 52852 71000 52910
rect 70802 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70802 52748 71000 52806
rect 70802 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70802 52644 71000 52702
rect 70802 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70802 52540 71000 52598
rect 70802 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70802 52436 71000 52494
rect 70802 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70802 52332 71000 52390
rect 70802 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70802 52228 71000 52286
rect 70802 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70802 52124 71000 52182
rect 70802 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70802 52020 71000 52078
rect 70802 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70802 51916 71000 51974
rect 70802 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70802 51812 71000 51870
rect 70802 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70802 51708 71000 51766
rect 70802 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70802 51604 71000 51662
rect 70802 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70802 51500 71000 51558
rect 70802 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70802 51396 71000 51454
rect 70802 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70802 51292 71000 51350
rect 70802 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70802 51188 71000 51246
rect 70802 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70802 51084 71000 51142
rect 70802 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70802 50980 71000 51038
rect 70802 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70802 50876 71000 50934
rect 70802 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70802 50772 71000 50830
rect 70802 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70802 50668 71000 50726
rect 70802 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70802 50564 71000 50622
rect 70802 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70802 50460 71000 50518
rect 70802 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70802 50356 71000 50414
rect 70802 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70802 50252 71000 50310
rect 70802 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70802 50148 71000 50206
rect 70802 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70802 50044 71000 50102
rect 70802 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70802 49940 71000 49998
rect 70802 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70802 49836 71000 49894
rect 70802 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70802 49732 71000 49790
rect 70802 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70802 49628 71000 49686
rect 70802 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70802 49524 71000 49582
rect 70802 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70802 49420 71000 49478
rect 70802 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70802 49316 71000 49374
rect 70802 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70802 49212 71000 49270
rect 70802 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70802 49108 71000 49166
rect 70802 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70802 49004 71000 49062
rect 70802 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70802 48900 71000 48958
rect 70802 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70802 48796 71000 48854
rect 70802 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70802 48692 71000 48750
rect 70802 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70802 48588 71000 48646
rect 70802 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70802 48484 71000 48542
rect 70802 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70802 48380 71000 48438
rect 70802 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70802 48276 71000 48334
rect 70802 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70802 48172 71000 48230
rect 70802 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70802 48068 71000 48126
rect 70802 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70802 47964 71000 48022
rect 70802 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70802 47860 71000 47918
rect 70802 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70802 47756 71000 47814
rect 70802 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70802 47652 71000 47710
rect 70802 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70802 47548 71000 47606
rect 70802 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70802 47444 71000 47502
rect 70802 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70802 47340 71000 47398
rect 70802 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70802 47236 71000 47294
rect 70802 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70802 47132 71000 47190
rect 70802 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70802 47028 71000 47086
rect 70802 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70802 46924 71000 46982
rect 70802 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70802 46820 71000 46878
rect 70802 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70802 46716 71000 46774
rect 70802 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70802 46612 71000 46670
rect 70802 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70802 46508 71000 46566
rect 70802 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70802 46404 71000 46462
rect 70802 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70802 46300 71000 46358
rect 70802 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70802 46196 71000 46254
rect 70802 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70802 46092 71000 46150
rect 70802 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70802 45988 71000 46046
rect 70802 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70802 45884 71000 45942
rect 70802 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70802 45780 71000 45838
rect 70802 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70802 45676 71000 45734
rect 70802 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70802 45572 71000 45630
rect 70802 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70802 45468 71000 45526
rect 70802 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70802 45364 71000 45422
rect 70802 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70802 45260 71000 45318
rect 70802 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70802 45156 71000 45214
rect 70802 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70802 45052 71000 45110
rect 70802 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70802 44948 71000 45006
tri 13291 44921 13295 44925 sw
rect 13097 44913 13295 44921
tri 13295 44913 13303 44921 sw
rect 13097 44905 13303 44913
tri 13303 44905 13311 44913 sw
rect 13097 44897 13311 44905
tri 13311 44897 13319 44905 sw
rect 70802 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13097 44889 13319 44897
tri 13319 44889 13327 44897 sw
rect 13097 44881 13327 44889
tri 13327 44881 13335 44889 sw
rect 13097 44877 13335 44881
tri 13335 44877 13339 44881 sw
rect 13097 44869 13339 44877
tri 13339 44869 13347 44877 sw
rect 13097 44861 13347 44869
tri 13347 44861 13355 44869 sw
rect 13097 44853 13355 44861
tri 13355 44853 13363 44861 sw
rect 13097 44845 13363 44853
tri 13363 44845 13371 44853 sw
rect 13097 44843 13371 44845
tri 13097 44839 13101 44843 ne
rect 13101 44839 13371 44843
tri 13101 44831 13109 44839 ne
rect 13109 44837 13371 44839
tri 13371 44837 13379 44845 sw
rect 70802 44844 71000 44902
rect 13109 44831 13379 44837
tri 13109 44823 13117 44831 ne
rect 13117 44829 13379 44831
tri 13379 44829 13387 44837 sw
rect 13117 44824 13387 44829
rect 13117 44823 13254 44824
tri 13117 44815 13125 44823 ne
rect 13125 44815 13254 44823
tri 13125 44807 13133 44815 ne
rect 13133 44807 13254 44815
tri 13133 44799 13141 44807 ne
rect 13141 44799 13254 44807
tri 13141 44791 13149 44799 ne
rect 13149 44791 13254 44799
tri 13149 44783 13157 44791 ne
rect 13157 44783 13254 44791
tri 13157 44775 13165 44783 ne
rect 13165 44778 13254 44783
rect 13300 44821 13387 44824
tri 13387 44821 13395 44829 sw
rect 13300 44813 13395 44821
tri 13395 44813 13403 44821 sw
rect 13300 44805 13403 44813
tri 13403 44805 13411 44813 sw
rect 13300 44797 13411 44805
tri 13411 44797 13419 44805 sw
rect 70802 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 13300 44789 13419 44797
tri 13419 44789 13427 44797 sw
rect 13300 44781 13427 44789
tri 13427 44781 13435 44789 sw
rect 13300 44778 13435 44781
rect 13165 44775 13435 44778
tri 13165 44772 13168 44775 ne
rect 13168 44773 13435 44775
tri 13435 44773 13443 44781 sw
rect 13168 44772 13443 44773
tri 13168 44764 13176 44772 ne
rect 13176 44765 13443 44772
tri 13443 44765 13451 44773 sw
rect 13176 44764 13451 44765
tri 13176 44756 13184 44764 ne
rect 13184 44757 13451 44764
tri 13451 44757 13459 44765 sw
rect 13184 44756 13459 44757
tri 13184 44748 13192 44756 ne
rect 13192 44749 13459 44756
tri 13459 44749 13467 44757 sw
rect 13192 44748 13467 44749
tri 13192 44740 13200 44748 ne
rect 13200 44743 13467 44748
tri 13467 44743 13473 44749 sw
rect 13200 44740 13473 44743
tri 13200 44732 13208 44740 ne
rect 13208 44735 13473 44740
tri 13473 44735 13481 44743 sw
rect 70802 44740 71000 44798
rect 13208 44732 13481 44735
tri 13208 44724 13216 44732 ne
rect 13216 44727 13481 44732
tri 13481 44727 13489 44735 sw
rect 13216 44724 13489 44727
tri 13216 44716 13224 44724 ne
rect 13224 44719 13489 44724
tri 13489 44719 13497 44727 sw
rect 13224 44716 13497 44719
tri 13224 44708 13232 44716 ne
rect 13232 44711 13497 44716
tri 13497 44711 13505 44719 sw
rect 13232 44708 13505 44711
tri 13232 44700 13240 44708 ne
rect 13240 44703 13505 44708
tri 13505 44703 13513 44711 sw
rect 13240 44700 13513 44703
tri 13240 44692 13248 44700 ne
rect 13248 44695 13513 44700
tri 13513 44695 13521 44703 sw
rect 13248 44692 13521 44695
tri 13248 44684 13256 44692 ne
rect 13256 44684 13386 44692
tri 13256 44679 13261 44684 ne
rect 13261 44679 13386 44684
tri 13261 44671 13269 44679 ne
rect 13269 44671 13386 44679
tri 13269 44663 13277 44671 ne
rect 13277 44663 13386 44671
tri 13277 44655 13285 44663 ne
rect 13285 44655 13386 44663
tri 13285 44647 13293 44655 ne
rect 13293 44647 13386 44655
tri 13293 44639 13301 44647 ne
rect 13301 44646 13386 44647
rect 13432 44687 13521 44692
tri 13521 44687 13529 44695 sw
rect 70802 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 13432 44679 13529 44687
tri 13529 44679 13537 44687 sw
rect 13432 44671 13537 44679
tri 13537 44671 13545 44679 sw
rect 13432 44663 13545 44671
tri 13545 44663 13553 44671 sw
rect 13432 44655 13553 44663
tri 13553 44655 13561 44663 sw
rect 13432 44647 13561 44655
tri 13561 44647 13569 44655 sw
rect 13432 44646 13569 44647
rect 13301 44639 13569 44646
tri 13569 44639 13577 44647 sw
tri 13301 44631 13309 44639 ne
rect 13309 44631 13577 44639
tri 13577 44631 13585 44639 sw
rect 70802 44636 71000 44694
tri 13309 44623 13317 44631 ne
rect 13317 44623 13585 44631
tri 13585 44623 13593 44631 sw
tri 13317 44615 13325 44623 ne
rect 13325 44615 13593 44623
tri 13593 44615 13601 44623 sw
tri 13325 44607 13333 44615 ne
rect 13333 44607 13601 44615
tri 13601 44607 13609 44615 sw
tri 13333 44601 13339 44607 ne
rect 13339 44601 13609 44607
tri 13609 44601 13615 44607 sw
tri 13339 44593 13347 44601 ne
rect 13347 44593 13615 44601
tri 13615 44593 13623 44601 sw
tri 13347 44585 13355 44593 ne
rect 13355 44585 13623 44593
tri 13623 44585 13631 44593 sw
rect 70802 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13355 44577 13363 44585 ne
rect 13363 44577 13631 44585
tri 13631 44577 13639 44585 sw
tri 13363 44569 13371 44577 ne
rect 13371 44569 13639 44577
tri 13639 44569 13647 44577 sw
tri 13371 44561 13379 44569 ne
rect 13379 44561 13647 44569
tri 13647 44561 13655 44569 sw
tri 13379 44553 13387 44561 ne
rect 13387 44560 13655 44561
rect 13387 44553 13518 44560
tri 13387 44545 13395 44553 ne
rect 13395 44545 13518 44553
tri 13395 44537 13403 44545 ne
rect 13403 44537 13518 44545
tri 13403 44529 13411 44537 ne
rect 13411 44529 13518 44537
tri 13411 44521 13419 44529 ne
rect 13419 44521 13518 44529
tri 13419 44513 13427 44521 ne
rect 13427 44514 13518 44521
rect 13564 44553 13655 44560
tri 13655 44553 13663 44561 sw
rect 13564 44545 13663 44553
tri 13663 44545 13671 44553 sw
rect 13564 44537 13671 44545
tri 13671 44537 13679 44545 sw
rect 13564 44529 13679 44537
tri 13679 44529 13687 44537 sw
rect 70802 44532 71000 44590
rect 13564 44521 13687 44529
tri 13687 44521 13695 44529 sw
rect 13564 44514 13695 44521
rect 13427 44513 13695 44514
tri 13695 44513 13703 44521 sw
tri 13427 44505 13435 44513 ne
rect 13435 44505 13703 44513
tri 13703 44505 13711 44513 sw
tri 13435 44497 13443 44505 ne
rect 13443 44497 13711 44505
tri 13711 44497 13719 44505 sw
tri 13443 44489 13451 44497 ne
rect 13451 44489 13719 44497
tri 13719 44489 13727 44497 sw
tri 13451 44481 13459 44489 ne
rect 13459 44481 13727 44489
tri 13727 44481 13735 44489 sw
rect 70802 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
tri 13459 44473 13467 44481 ne
rect 13467 44473 13735 44481
tri 13735 44473 13743 44481 sw
tri 13467 44465 13475 44473 ne
rect 13475 44465 13743 44473
tri 13743 44465 13751 44473 sw
tri 13475 44459 13481 44465 ne
rect 13481 44459 13751 44465
tri 13751 44459 13757 44465 sw
tri 13481 44451 13489 44459 ne
rect 13489 44451 13757 44459
tri 13757 44451 13765 44459 sw
tri 13489 44443 13497 44451 ne
rect 13497 44443 13765 44451
tri 13765 44443 13773 44451 sw
tri 13497 44435 13505 44443 ne
rect 13505 44435 13773 44443
tri 13773 44435 13781 44443 sw
tri 13505 44427 13513 44435 ne
rect 13513 44428 13781 44435
rect 13513 44427 13650 44428
tri 13513 44419 13521 44427 ne
rect 13521 44419 13650 44427
tri 13521 44411 13529 44419 ne
rect 13529 44411 13650 44419
tri 13529 44403 13537 44411 ne
rect 13537 44403 13650 44411
tri 13537 44395 13545 44403 ne
rect 13545 44395 13650 44403
tri 13545 44387 13553 44395 ne
rect 13553 44387 13650 44395
tri 13553 44379 13561 44387 ne
rect 13561 44382 13650 44387
rect 13696 44427 13781 44428
tri 13781 44427 13789 44435 sw
rect 70802 44428 71000 44486
rect 13696 44419 13789 44427
tri 13789 44419 13797 44427 sw
rect 13696 44411 13797 44419
tri 13797 44411 13805 44419 sw
rect 13696 44403 13805 44411
tri 13805 44403 13813 44411 sw
rect 13696 44395 13813 44403
tri 13813 44395 13821 44403 sw
rect 13696 44387 13821 44395
tri 13821 44387 13829 44395 sw
rect 13696 44382 13829 44387
rect 13561 44379 13829 44382
tri 13829 44379 13837 44387 sw
rect 70802 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
tri 13561 44371 13569 44379 ne
rect 13569 44371 13837 44379
tri 13837 44371 13845 44379 sw
tri 13569 44363 13577 44371 ne
rect 13577 44363 13845 44371
tri 13845 44363 13853 44371 sw
tri 13577 44355 13585 44363 ne
rect 13585 44355 13853 44363
tri 13853 44355 13861 44363 sw
tri 13585 44347 13593 44355 ne
rect 13593 44347 13861 44355
tri 13861 44347 13869 44355 sw
tri 13593 44339 13601 44347 ne
rect 13601 44346 13869 44347
tri 13869 44346 13870 44347 sw
rect 13601 44339 13870 44346
tri 13601 44331 13609 44339 ne
rect 13609 44338 13870 44339
tri 13870 44338 13878 44346 sw
rect 13609 44331 13878 44338
tri 13609 44323 13617 44331 ne
rect 13617 44330 13878 44331
tri 13878 44330 13886 44338 sw
rect 13617 44323 13886 44330
tri 13617 44322 13618 44323 ne
rect 13618 44322 13886 44323
tri 13886 44322 13894 44330 sw
rect 70802 44324 71000 44382
tri 13618 44314 13626 44322 ne
rect 13626 44314 13894 44322
tri 13894 44314 13902 44322 sw
tri 13626 44306 13634 44314 ne
rect 13634 44306 13902 44314
tri 13902 44306 13910 44314 sw
tri 13634 44298 13642 44306 ne
rect 13642 44298 13910 44306
tri 13910 44298 13918 44306 sw
tri 13642 44290 13650 44298 ne
rect 13650 44296 13918 44298
rect 13650 44290 13782 44296
tri 13650 44282 13658 44290 ne
rect 13658 44282 13782 44290
tri 13658 44274 13666 44282 ne
rect 13666 44274 13782 44282
tri 13666 44266 13674 44274 ne
rect 13674 44266 13782 44274
tri 13674 44258 13682 44266 ne
rect 13682 44258 13782 44266
tri 13682 44250 13690 44258 ne
rect 13690 44250 13782 44258
rect 13828 44290 13918 44296
tri 13918 44290 13926 44298 sw
rect 13828 44282 13926 44290
tri 13926 44282 13934 44290 sw
rect 13828 44274 13934 44282
tri 13934 44274 13942 44282 sw
rect 70802 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 13828 44266 13942 44274
tri 13942 44266 13950 44274 sw
rect 13828 44258 13950 44266
tri 13950 44258 13958 44266 sw
rect 13828 44255 13958 44258
tri 13958 44255 13961 44258 sw
rect 13828 44250 13961 44255
tri 13690 44242 13698 44250 ne
rect 13698 44247 13961 44250
tri 13961 44247 13969 44255 sw
rect 13698 44242 13969 44247
tri 13698 44234 13706 44242 ne
rect 13706 44239 13969 44242
tri 13969 44239 13977 44247 sw
rect 13706 44234 13977 44239
tri 13706 44226 13714 44234 ne
rect 13714 44231 13977 44234
tri 13977 44231 13985 44239 sw
rect 13714 44226 13985 44231
tri 13714 44218 13722 44226 ne
rect 13722 44223 13985 44226
tri 13985 44223 13993 44231 sw
rect 13722 44218 13993 44223
tri 13722 44215 13725 44218 ne
rect 13725 44215 13993 44218
tri 13993 44215 14001 44223 sw
rect 70802 44220 71000 44278
tri 13725 44207 13733 44215 ne
rect 13733 44207 14001 44215
tri 14001 44207 14009 44215 sw
tri 13733 44199 13741 44207 ne
rect 13741 44199 14009 44207
tri 14009 44199 14017 44207 sw
tri 13741 44191 13749 44199 ne
rect 13749 44191 14017 44199
tri 14017 44191 14025 44199 sw
tri 13749 44183 13757 44191 ne
rect 13757 44183 14025 44191
tri 14025 44183 14033 44191 sw
tri 13757 44175 13765 44183 ne
rect 13765 44175 14033 44183
tri 14033 44175 14041 44183 sw
tri 13765 44167 13773 44175 ne
rect 13773 44167 14041 44175
tri 14041 44167 14049 44175 sw
rect 70802 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
tri 13773 44159 13781 44167 ne
rect 13781 44164 14049 44167
rect 13781 44159 13914 44164
tri 13781 44151 13789 44159 ne
rect 13789 44151 13914 44159
tri 13789 44143 13797 44151 ne
rect 13797 44143 13914 44151
tri 13797 44135 13805 44143 ne
rect 13805 44135 13914 44143
tri 13805 44127 13813 44135 ne
rect 13813 44127 13914 44135
tri 13813 44119 13821 44127 ne
rect 13821 44119 13914 44127
tri 13821 44111 13829 44119 ne
rect 13829 44118 13914 44119
rect 13960 44159 14049 44164
tri 14049 44159 14057 44167 sw
rect 13960 44151 14057 44159
tri 14057 44151 14065 44159 sw
rect 13960 44143 14065 44151
tri 14065 44143 14073 44151 sw
rect 13960 44135 14073 44143
tri 14073 44135 14081 44143 sw
rect 13960 44127 14081 44135
tri 14081 44127 14089 44135 sw
rect 13960 44119 14089 44127
tri 14089 44119 14097 44127 sw
rect 13960 44118 14097 44119
rect 13829 44111 14097 44118
tri 14097 44111 14105 44119 sw
rect 70802 44116 71000 44174
tri 13829 44103 13837 44111 ne
rect 13837 44103 14105 44111
tri 14105 44103 14113 44111 sw
tri 13837 44101 13839 44103 ne
rect 13839 44101 14113 44103
tri 13839 44093 13847 44101 ne
rect 13847 44095 14113 44101
tri 14113 44095 14121 44103 sw
rect 13847 44093 14121 44095
tri 13847 44085 13855 44093 ne
rect 13855 44087 14121 44093
tri 14121 44087 14129 44095 sw
rect 13855 44085 14129 44087
tri 13855 44077 13863 44085 ne
rect 13863 44079 14129 44085
tri 14129 44079 14137 44087 sw
rect 13863 44077 14137 44079
tri 13863 44069 13871 44077 ne
rect 13871 44071 14137 44077
tri 14137 44071 14145 44079 sw
rect 13871 44069 14145 44071
tri 13871 44061 13879 44069 ne
rect 13879 44063 14145 44069
tri 14145 44063 14153 44071 sw
rect 70802 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 13879 44061 14153 44063
tri 13879 44053 13887 44061 ne
rect 13887 44055 14153 44061
tri 14153 44055 14161 44063 sw
rect 13887 44053 14161 44055
tri 13887 44045 13895 44053 ne
rect 13895 44047 14161 44053
tri 14161 44047 14169 44055 sw
rect 13895 44045 14169 44047
tri 13895 44037 13903 44045 ne
rect 13903 44039 14169 44045
tri 14169 44039 14177 44047 sw
rect 13903 44037 14177 44039
tri 13903 44029 13911 44037 ne
rect 13911 44032 14177 44037
rect 13911 44029 14046 44032
tri 13911 44021 13919 44029 ne
rect 13919 44021 14046 44029
tri 13919 44013 13927 44021 ne
rect 13927 44013 14046 44021
tri 13927 44005 13935 44013 ne
rect 13935 44005 14046 44013
tri 13935 43997 13943 44005 ne
rect 13943 43997 14046 44005
tri 13943 43991 13949 43997 ne
rect 13949 43991 14046 43997
tri 13949 43983 13957 43991 ne
rect 13957 43986 14046 43991
rect 14092 44031 14177 44032
tri 14177 44031 14185 44039 sw
rect 14092 44023 14185 44031
tri 14185 44023 14193 44031 sw
rect 14092 44015 14193 44023
tri 14193 44015 14201 44023 sw
rect 14092 44007 14201 44015
tri 14201 44007 14209 44015 sw
rect 70802 44012 71000 44070
rect 14092 43999 14209 44007
tri 14209 43999 14217 44007 sw
rect 14092 43991 14217 43999
tri 14217 43991 14225 43999 sw
rect 14092 43986 14225 43991
rect 13957 43983 14225 43986
tri 14225 43983 14233 43991 sw
tri 13957 43975 13965 43983 ne
rect 13965 43975 14233 43983
tri 14233 43975 14241 43983 sw
tri 13965 43967 13973 43975 ne
rect 13973 43967 14241 43975
tri 14241 43967 14249 43975 sw
tri 13973 43959 13981 43967 ne
rect 13981 43959 14249 43967
tri 14249 43959 14257 43967 sw
rect 70802 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13981 43951 13989 43959 ne
rect 13989 43951 14257 43959
tri 14257 43951 14265 43959 sw
tri 13989 43943 13997 43951 ne
rect 13997 43943 14265 43951
tri 14265 43943 14273 43951 sw
tri 13997 43935 14005 43943 ne
rect 14005 43935 14273 43943
tri 14273 43935 14281 43943 sw
tri 14005 43927 14013 43935 ne
rect 14013 43927 14281 43935
tri 14281 43927 14289 43935 sw
tri 14013 43919 14021 43927 ne
rect 14021 43919 14289 43927
tri 14289 43919 14297 43927 sw
tri 14021 43911 14029 43919 ne
rect 14029 43911 14297 43919
tri 14297 43911 14305 43919 sw
tri 14029 43903 14037 43911 ne
rect 14037 43903 14305 43911
tri 14305 43903 14313 43911 sw
rect 70802 43908 71000 43966
tri 14037 43895 14045 43903 ne
rect 14045 43900 14313 43903
rect 14045 43895 14178 43900
tri 14045 43887 14053 43895 ne
rect 14053 43887 14178 43895
tri 14053 43883 14057 43887 ne
rect 14057 43883 14178 43887
tri 14057 43875 14065 43883 ne
rect 14065 43875 14178 43883
tri 14065 43867 14073 43875 ne
rect 14073 43867 14178 43875
tri 14073 43859 14081 43867 ne
rect 14081 43859 14178 43867
tri 14081 43851 14089 43859 ne
rect 14089 43854 14178 43859
rect 14224 43895 14313 43900
tri 14313 43895 14321 43903 sw
rect 14224 43887 14321 43895
tri 14321 43887 14329 43895 sw
rect 14224 43883 14329 43887
tri 14329 43883 14333 43887 sw
rect 14224 43875 14333 43883
tri 14333 43875 14341 43883 sw
rect 14224 43867 14341 43875
tri 14341 43867 14349 43875 sw
rect 14224 43859 14349 43867
tri 14349 43859 14357 43867 sw
rect 70802 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 14224 43854 14357 43859
rect 14089 43851 14357 43854
tri 14357 43851 14365 43859 sw
tri 14089 43843 14097 43851 ne
rect 14097 43843 14365 43851
tri 14365 43843 14373 43851 sw
tri 14097 43835 14105 43843 ne
rect 14105 43835 14373 43843
tri 14373 43835 14381 43843 sw
tri 14105 43827 14113 43835 ne
rect 14113 43827 14381 43835
tri 14381 43827 14389 43835 sw
tri 14113 43819 14121 43827 ne
rect 14121 43825 14389 43827
tri 14389 43825 14391 43827 sw
rect 14121 43819 14391 43825
tri 14121 43811 14129 43819 ne
rect 14129 43817 14391 43819
tri 14391 43817 14399 43825 sw
rect 14129 43811 14399 43817
tri 14129 43803 14137 43811 ne
rect 14137 43809 14399 43811
tri 14399 43809 14407 43817 sw
rect 14137 43803 14407 43809
tri 14137 43795 14145 43803 ne
rect 14145 43801 14407 43803
tri 14407 43801 14415 43809 sw
rect 70802 43804 71000 43862
rect 14145 43795 14415 43801
tri 14145 43787 14153 43795 ne
rect 14153 43793 14415 43795
tri 14415 43793 14423 43801 sw
rect 14153 43787 14423 43793
tri 14153 43779 14161 43787 ne
rect 14161 43785 14423 43787
tri 14423 43785 14431 43793 sw
rect 14161 43779 14431 43785
tri 14161 43771 14169 43779 ne
rect 14169 43777 14431 43779
tri 14431 43777 14439 43785 sw
rect 14169 43771 14439 43777
tri 14169 43763 14177 43771 ne
rect 14177 43769 14439 43771
tri 14439 43769 14447 43777 sw
rect 14177 43768 14447 43769
rect 14177 43763 14310 43768
tri 14177 43755 14185 43763 ne
rect 14185 43755 14310 43763
tri 14185 43747 14193 43755 ne
rect 14193 43747 14310 43755
tri 14193 43742 14198 43747 ne
rect 14198 43742 14310 43747
tri 14198 43734 14206 43742 ne
rect 14206 43734 14310 43742
tri 14206 43726 14214 43734 ne
rect 14214 43726 14310 43734
tri 14214 43718 14222 43726 ne
rect 14222 43722 14310 43726
rect 14356 43761 14447 43768
tri 14447 43761 14455 43769 sw
rect 14356 43753 14455 43761
tri 14455 43753 14463 43761 sw
rect 70802 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43745 14463 43753
tri 14463 43745 14471 43753 sw
rect 14356 43737 14471 43745
tri 14471 43737 14479 43745 sw
rect 14356 43729 14479 43737
tri 14479 43729 14487 43737 sw
rect 14356 43723 14487 43729
tri 14487 43723 14493 43729 sw
rect 14356 43722 14493 43723
rect 14222 43718 14493 43722
tri 14222 43710 14230 43718 ne
rect 14230 43715 14493 43718
tri 14493 43715 14501 43723 sw
rect 14230 43710 14501 43715
tri 14230 43702 14238 43710 ne
rect 14238 43707 14501 43710
tri 14501 43707 14509 43715 sw
rect 14238 43702 14509 43707
tri 14238 43694 14246 43702 ne
rect 14246 43699 14509 43702
tri 14509 43699 14517 43707 sw
rect 70802 43700 71000 43758
rect 14246 43694 14517 43699
tri 14246 43686 14254 43694 ne
rect 14254 43691 14517 43694
tri 14517 43691 14525 43699 sw
rect 14254 43686 14525 43691
tri 14254 43678 14262 43686 ne
rect 14262 43683 14525 43686
tri 14525 43683 14533 43691 sw
rect 14262 43678 14533 43683
tri 14262 43670 14270 43678 ne
rect 14270 43675 14533 43678
tri 14533 43675 14541 43683 sw
rect 14270 43670 14541 43675
tri 14270 43662 14278 43670 ne
rect 14278 43667 14541 43670
tri 14541 43667 14549 43675 sw
rect 14278 43662 14549 43667
tri 14278 43654 14286 43662 ne
rect 14286 43659 14549 43662
tri 14549 43659 14557 43667 sw
rect 14286 43654 14557 43659
tri 14286 43646 14294 43654 ne
rect 14294 43651 14557 43654
tri 14557 43651 14565 43659 sw
rect 70802 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14294 43646 14565 43651
tri 14294 43638 14302 43646 ne
rect 14302 43643 14565 43646
tri 14565 43643 14573 43651 sw
rect 14302 43638 14573 43643
tri 14302 43630 14310 43638 ne
rect 14310 43636 14573 43638
rect 14310 43630 14442 43636
tri 14310 43622 14318 43630 ne
rect 14318 43622 14442 43630
tri 14318 43614 14326 43622 ne
rect 14326 43614 14442 43622
tri 14326 43606 14334 43614 ne
rect 14334 43606 14442 43614
tri 14334 43599 14341 43606 ne
rect 14341 43599 14442 43606
tri 14341 43591 14349 43599 ne
rect 14349 43591 14442 43599
tri 14349 43583 14357 43591 ne
rect 14357 43590 14442 43591
rect 14488 43635 14573 43636
tri 14573 43635 14581 43643 sw
rect 14488 43627 14581 43635
tri 14581 43627 14589 43635 sw
rect 14488 43619 14589 43627
tri 14589 43619 14597 43627 sw
rect 14488 43611 14597 43619
tri 14597 43611 14605 43619 sw
rect 14488 43603 14605 43611
tri 14605 43603 14613 43611 sw
rect 14488 43599 14613 43603
tri 14613 43599 14617 43603 sw
rect 14488 43591 14617 43599
tri 14617 43591 14625 43599 sw
rect 70802 43596 71000 43654
rect 14488 43590 14625 43591
rect 14357 43583 14625 43590
tri 14625 43583 14633 43591 sw
tri 14357 43575 14365 43583 ne
rect 14365 43575 14633 43583
tri 14633 43575 14641 43583 sw
tri 14365 43567 14373 43575 ne
rect 14373 43567 14641 43575
tri 14641 43567 14649 43575 sw
tri 14373 43559 14381 43567 ne
rect 14381 43559 14649 43567
tri 14649 43559 14657 43567 sw
tri 14381 43556 14384 43559 ne
rect 14384 43556 14657 43559
tri 14384 43551 14389 43556 ne
rect 14389 43551 14657 43556
tri 14657 43551 14665 43559 sw
tri 14389 43543 14397 43551 ne
rect 14397 43543 14665 43551
tri 14665 43543 14673 43551 sw
rect 70802 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
tri 14397 43535 14405 43543 ne
rect 14405 43535 14673 43543
tri 14673 43535 14681 43543 sw
tri 14405 43527 14413 43535 ne
rect 14413 43527 14681 43535
tri 14681 43527 14689 43535 sw
tri 14413 43519 14421 43527 ne
rect 14421 43519 14689 43527
tri 14689 43519 14697 43527 sw
tri 14421 43511 14429 43519 ne
rect 14429 43511 14697 43519
tri 14697 43511 14705 43519 sw
tri 14429 43503 14437 43511 ne
rect 14437 43504 14705 43511
rect 14437 43503 14574 43504
tri 14437 43495 14445 43503 ne
rect 14445 43495 14574 43503
tri 14445 43487 14453 43495 ne
rect 14453 43487 14574 43495
tri 14453 43479 14461 43487 ne
rect 14461 43479 14574 43487
tri 14461 43471 14469 43479 ne
rect 14469 43471 14574 43479
tri 14469 43470 14470 43471 ne
rect 14470 43470 14574 43471
tri 14470 43462 14478 43470 ne
rect 14478 43462 14574 43470
tri 14478 43454 14486 43462 ne
rect 14486 43458 14574 43462
rect 14620 43503 14705 43504
tri 14705 43503 14713 43511 sw
rect 14620 43495 14713 43503
tri 14713 43495 14721 43503 sw
rect 14620 43487 14721 43495
tri 14721 43487 14729 43495 sw
rect 70802 43492 71000 43550
rect 14620 43479 14729 43487
tri 14729 43479 14737 43487 sw
rect 14620 43471 14737 43479
tri 14737 43471 14745 43479 sw
rect 14620 43470 14745 43471
tri 14745 43470 14746 43471 sw
rect 14620 43462 14746 43470
tri 14746 43462 14754 43470 sw
rect 14620 43458 14754 43462
rect 14486 43454 14754 43458
tri 14754 43454 14762 43462 sw
tri 14486 43446 14494 43454 ne
rect 14494 43446 14762 43454
tri 14762 43446 14770 43454 sw
rect 70802 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14494 43438 14502 43446 ne
rect 14502 43438 14770 43446
tri 14770 43438 14778 43446 sw
tri 14502 43430 14510 43438 ne
rect 14510 43430 14778 43438
tri 14778 43430 14786 43438 sw
tri 14510 43422 14518 43430 ne
rect 14518 43422 14786 43430
tri 14786 43422 14794 43430 sw
tri 14518 43414 14526 43422 ne
rect 14526 43414 14794 43422
tri 14794 43414 14802 43422 sw
tri 14526 43406 14534 43414 ne
rect 14534 43406 14802 43414
tri 14802 43406 14810 43414 sw
tri 14534 43398 14542 43406 ne
rect 14542 43398 14810 43406
tri 14810 43398 14818 43406 sw
tri 14542 43390 14550 43398 ne
rect 14550 43390 14818 43398
tri 14818 43390 14826 43398 sw
tri 14550 43382 14558 43390 ne
rect 14558 43382 14826 43390
tri 14826 43382 14834 43390 sw
rect 70802 43388 71000 43446
tri 14558 43374 14566 43382 ne
rect 14566 43374 14834 43382
tri 14834 43374 14842 43382 sw
tri 14566 43366 14574 43374 ne
rect 14574 43372 14842 43374
rect 14574 43366 14706 43372
tri 14574 43358 14582 43366 ne
rect 14582 43358 14706 43366
tri 14582 43350 14590 43358 ne
rect 14590 43350 14706 43358
tri 14590 43342 14598 43350 ne
rect 14598 43342 14706 43350
tri 14598 43339 14601 43342 ne
rect 14601 43339 14706 43342
tri 14601 43331 14609 43339 ne
rect 14609 43331 14706 43339
tri 14609 43323 14617 43331 ne
rect 14617 43326 14706 43331
rect 14752 43366 14842 43372
tri 14842 43366 14850 43374 sw
rect 14752 43358 14850 43366
tri 14850 43358 14858 43366 sw
rect 14752 43350 14858 43358
tri 14858 43350 14866 43358 sw
rect 14752 43342 14866 43350
tri 14866 43342 14874 43350 sw
rect 70802 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 14752 43339 14874 43342
tri 14874 43339 14877 43342 sw
rect 14752 43331 14877 43339
tri 14877 43331 14885 43339 sw
rect 14752 43326 14885 43331
rect 14617 43323 14885 43326
tri 14885 43323 14893 43331 sw
tri 14617 43315 14625 43323 ne
rect 14625 43315 14893 43323
tri 14893 43315 14901 43323 sw
tri 14625 43307 14633 43315 ne
rect 14633 43307 14901 43315
tri 14901 43307 14909 43315 sw
tri 14633 43299 14641 43307 ne
rect 14641 43299 14909 43307
tri 14909 43299 14917 43307 sw
tri 14641 43291 14649 43299 ne
rect 14649 43291 14917 43299
tri 14917 43291 14925 43299 sw
tri 14649 43283 14657 43291 ne
rect 14657 43283 14925 43291
tri 14925 43283 14933 43291 sw
rect 70802 43284 71000 43342
tri 14657 43275 14665 43283 ne
rect 14665 43275 14933 43283
tri 14933 43275 14941 43283 sw
tri 14665 43267 14673 43275 ne
rect 14673 43267 14941 43275
tri 14941 43267 14949 43275 sw
tri 14673 43259 14681 43267 ne
rect 14681 43259 14949 43267
tri 14949 43259 14957 43267 sw
tri 14681 43251 14689 43259 ne
rect 14689 43251 14957 43259
tri 14957 43251 14965 43259 sw
tri 14689 43243 14697 43251 ne
rect 14697 43243 14965 43251
tri 14965 43243 14973 43251 sw
tri 14697 43235 14705 43243 ne
rect 14705 43240 14973 43243
rect 14705 43235 14838 43240
tri 14705 43227 14713 43235 ne
rect 14713 43227 14838 43235
tri 14713 43219 14721 43227 ne
rect 14721 43219 14838 43227
tri 14721 43211 14729 43219 ne
rect 14729 43211 14838 43219
tri 14729 43203 14737 43211 ne
rect 14737 43203 14838 43211
tri 14737 43195 14745 43203 ne
rect 14745 43195 14838 43203
tri 14745 43194 14746 43195 ne
rect 14746 43194 14838 43195
rect 14884 43235 14973 43240
tri 14973 43235 14981 43243 sw
rect 70802 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43227 14981 43235
tri 14981 43227 14989 43235 sw
rect 14884 43219 14989 43227
tri 14989 43219 14997 43227 sw
rect 14884 43211 14997 43219
tri 14997 43211 15005 43219 sw
rect 14884 43203 15005 43211
tri 15005 43203 15013 43211 sw
rect 14884 43195 15013 43203
tri 15013 43195 15021 43203 sw
rect 14884 43194 15021 43195
tri 15021 43194 15022 43195 sw
tri 14746 43186 14754 43194 ne
rect 14754 43186 15022 43194
tri 15022 43186 15030 43194 sw
tri 14754 43178 14762 43186 ne
rect 14762 43178 15030 43186
tri 15030 43178 15038 43186 sw
rect 70802 43180 71000 43238
tri 14762 43170 14770 43178 ne
rect 14770 43170 15038 43178
tri 15038 43170 15046 43178 sw
tri 14770 43162 14778 43170 ne
rect 14778 43162 15046 43170
tri 15046 43162 15054 43170 sw
tri 14778 43154 14786 43162 ne
rect 14786 43154 15054 43162
tri 15054 43154 15062 43162 sw
tri 14786 43146 14794 43154 ne
rect 14794 43146 15062 43154
tri 15062 43146 15070 43154 sw
tri 14794 43138 14802 43146 ne
rect 14802 43138 15070 43146
tri 15070 43138 15078 43146 sw
tri 14802 43130 14810 43138 ne
rect 14810 43130 15078 43138
tri 15078 43130 15086 43138 sw
rect 70802 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14810 43122 14818 43130 ne
rect 14818 43122 15086 43130
tri 15086 43122 15094 43130 sw
tri 14818 43114 14826 43122 ne
rect 14826 43114 15094 43122
tri 15094 43114 15102 43122 sw
tri 14826 43106 14834 43114 ne
rect 14834 43108 15102 43114
rect 14834 43106 14970 43108
tri 14834 43098 14842 43106 ne
rect 14842 43098 14970 43106
tri 14842 43090 14850 43098 ne
rect 14850 43090 14970 43098
tri 14850 43082 14858 43090 ne
rect 14858 43082 14970 43090
tri 14858 43074 14866 43082 ne
rect 14866 43074 14970 43082
tri 14866 43066 14874 43074 ne
rect 14874 43066 14970 43074
tri 14874 43058 14882 43066 ne
rect 14882 43062 14970 43066
rect 15016 43106 15102 43108
tri 15102 43106 15110 43114 sw
rect 15016 43098 15110 43106
tri 15110 43098 15118 43106 sw
rect 15016 43090 15118 43098
tri 15118 43090 15126 43098 sw
rect 15016 43082 15126 43090
tri 15126 43082 15134 43090 sw
rect 15016 43074 15134 43082
tri 15134 43074 15142 43082 sw
rect 70802 43076 71000 43134
rect 15016 43066 15142 43074
tri 15142 43066 15150 43074 sw
rect 15016 43062 15150 43066
rect 14882 43058 15150 43062
tri 15150 43058 15158 43066 sw
tri 14882 43055 14885 43058 ne
rect 14885 43055 15158 43058
tri 15158 43055 15161 43058 sw
tri 14885 43047 14893 43055 ne
rect 14893 43047 15161 43055
tri 15161 43047 15169 43055 sw
tri 14893 43039 14901 43047 ne
rect 14901 43039 15169 43047
tri 15169 43039 15177 43047 sw
tri 14901 43031 14909 43039 ne
rect 14909 43031 15177 43039
tri 15177 43031 15185 43039 sw
tri 14909 43023 14917 43031 ne
rect 14917 43023 15185 43031
tri 15185 43023 15193 43031 sw
rect 70802 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14917 43015 14925 43023 ne
rect 14925 43015 15193 43023
tri 15193 43015 15201 43023 sw
tri 14925 43007 14933 43015 ne
rect 14933 43007 15201 43015
tri 15201 43007 15209 43015 sw
tri 14933 42999 14941 43007 ne
rect 14941 42999 15209 43007
tri 15209 42999 15217 43007 sw
tri 14941 42991 14949 42999 ne
rect 14949 42991 15217 42999
tri 15217 42991 15225 42999 sw
tri 14949 42983 14957 42991 ne
rect 14957 42983 15225 42991
tri 15225 42983 15233 42991 sw
tri 14957 42975 14965 42983 ne
rect 14965 42976 15233 42983
rect 14965 42975 15102 42976
tri 14965 42967 14973 42975 ne
rect 14973 42967 15102 42975
tri 14973 42959 14981 42967 ne
rect 14981 42959 15102 42967
tri 14981 42951 14989 42959 ne
rect 14989 42951 15102 42959
tri 14989 42943 14997 42951 ne
rect 14997 42943 15102 42951
tri 14997 42935 15005 42943 ne
rect 15005 42935 15102 42943
tri 15005 42927 15013 42935 ne
rect 15013 42930 15102 42935
rect 15148 42975 15233 42976
tri 15233 42975 15241 42983 sw
rect 15148 42967 15241 42975
tri 15241 42967 15249 42975 sw
rect 70802 42972 71000 43030
rect 15148 42959 15249 42967
tri 15249 42959 15257 42967 sw
rect 15148 42951 15257 42959
tri 15257 42951 15265 42959 sw
rect 15148 42943 15265 42951
tri 15265 42943 15273 42951 sw
rect 15148 42935 15273 42943
tri 15273 42935 15281 42943 sw
rect 15148 42930 15281 42935
rect 15013 42927 15281 42930
tri 15281 42927 15289 42935 sw
tri 15013 42924 15016 42927 ne
rect 15016 42924 15289 42927
tri 15289 42924 15292 42927 sw
rect 70802 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15016 42916 15024 42924 ne
rect 15024 42916 15292 42924
tri 15292 42916 15300 42924 sw
tri 15024 42908 15032 42916 ne
rect 15032 42908 15300 42916
tri 15300 42908 15308 42916 sw
tri 15032 42900 15040 42908 ne
rect 15040 42900 15308 42908
tri 15308 42900 15316 42908 sw
tri 15040 42892 15048 42900 ne
rect 15048 42892 15316 42900
tri 15316 42892 15324 42900 sw
tri 15048 42884 15056 42892 ne
rect 15056 42884 15324 42892
tri 15324 42884 15332 42892 sw
tri 15056 42876 15064 42884 ne
rect 15064 42876 15332 42884
tri 15332 42876 15340 42884 sw
tri 15064 42868 15072 42876 ne
rect 15072 42868 15340 42876
tri 15340 42868 15348 42876 sw
rect 70802 42868 71000 42926
tri 15072 42860 15080 42868 ne
rect 15080 42860 15348 42868
tri 15348 42860 15356 42868 sw
tri 15080 42852 15088 42860 ne
rect 15088 42852 15356 42860
tri 15356 42852 15364 42860 sw
tri 15088 42844 15096 42852 ne
rect 15096 42844 15364 42852
tri 15364 42844 15372 42852 sw
tri 15096 42836 15104 42844 ne
rect 15104 42836 15234 42844
tri 15104 42828 15112 42836 ne
rect 15112 42828 15234 42836
tri 15112 42820 15120 42828 ne
rect 15120 42820 15234 42828
tri 15120 42812 15128 42820 ne
rect 15128 42812 15234 42820
tri 15128 42804 15136 42812 ne
rect 15136 42804 15234 42812
tri 15136 42796 15144 42804 ne
rect 15144 42798 15234 42804
rect 15280 42836 15372 42844
tri 15372 42836 15380 42844 sw
rect 15280 42828 15380 42836
tri 15380 42828 15388 42836 sw
rect 15280 42820 15388 42828
tri 15388 42820 15396 42828 sw
rect 70802 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 15280 42812 15396 42820
tri 15396 42812 15404 42820 sw
rect 15280 42804 15404 42812
tri 15404 42804 15412 42812 sw
rect 15280 42798 15412 42804
rect 15144 42796 15412 42798
tri 15412 42796 15420 42804 sw
tri 15144 42788 15152 42796 ne
rect 15152 42788 15420 42796
tri 15420 42788 15428 42796 sw
tri 15152 42780 15160 42788 ne
rect 15160 42780 15428 42788
tri 15428 42780 15436 42788 sw
tri 15160 42779 15161 42780 ne
rect 15161 42779 15436 42780
tri 15436 42779 15437 42780 sw
tri 15161 42771 15169 42779 ne
rect 15169 42771 15437 42779
tri 15437 42771 15445 42779 sw
tri 15169 42763 15177 42771 ne
rect 15177 42763 15445 42771
tri 15445 42763 15453 42771 sw
rect 70802 42764 71000 42822
tri 15177 42755 15185 42763 ne
rect 15185 42755 15453 42763
tri 15453 42755 15461 42763 sw
tri 15185 42747 15193 42755 ne
rect 15193 42747 15461 42755
tri 15461 42747 15469 42755 sw
tri 15193 42739 15201 42747 ne
rect 15201 42739 15469 42747
tri 15469 42739 15477 42747 sw
tri 15201 42731 15209 42739 ne
rect 15209 42731 15477 42739
tri 15477 42731 15485 42739 sw
tri 15209 42723 15217 42731 ne
rect 15217 42723 15485 42731
tri 15485 42723 15493 42731 sw
tri 15217 42715 15225 42723 ne
rect 15225 42715 15493 42723
tri 15493 42715 15501 42723 sw
rect 70802 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
tri 15225 42707 15233 42715 ne
rect 15233 42712 15501 42715
rect 15233 42707 15366 42712
tri 15233 42699 15241 42707 ne
rect 15241 42699 15366 42707
tri 15241 42691 15249 42699 ne
rect 15249 42691 15366 42699
tri 15249 42683 15257 42691 ne
rect 15257 42683 15366 42691
tri 15257 42675 15265 42683 ne
rect 15265 42675 15366 42683
tri 15265 42667 15273 42675 ne
rect 15273 42667 15366 42675
tri 15273 42659 15281 42667 ne
rect 15281 42666 15366 42667
rect 15412 42707 15501 42712
tri 15501 42707 15509 42715 sw
rect 15412 42699 15509 42707
tri 15509 42699 15517 42707 sw
rect 15412 42691 15517 42699
tri 15517 42691 15525 42699 sw
rect 15412 42683 15525 42691
tri 15525 42683 15533 42691 sw
rect 15412 42675 15533 42683
tri 15533 42675 15541 42683 sw
rect 15412 42667 15541 42675
tri 15541 42667 15549 42675 sw
rect 15412 42666 15549 42667
rect 15281 42659 15549 42666
tri 15549 42659 15557 42667 sw
rect 70802 42660 71000 42718
tri 15281 42651 15289 42659 ne
rect 15289 42651 15557 42659
tri 15557 42651 15565 42659 sw
tri 15289 42643 15297 42651 ne
rect 15297 42643 15565 42651
tri 15565 42643 15573 42651 sw
tri 15297 42640 15300 42643 ne
rect 15300 42640 15573 42643
tri 15573 42640 15576 42643 sw
tri 15300 42632 15308 42640 ne
rect 15308 42632 15576 42640
tri 15576 42632 15584 42640 sw
tri 15308 42624 15316 42632 ne
rect 15316 42624 15584 42632
tri 15584 42624 15592 42632 sw
tri 15316 42616 15324 42624 ne
rect 15324 42616 15592 42624
tri 15592 42616 15600 42624 sw
tri 15324 42608 15332 42616 ne
rect 15332 42608 15600 42616
tri 15600 42608 15608 42616 sw
rect 70802 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15332 42600 15340 42608 ne
rect 15340 42600 15608 42608
tri 15608 42600 15616 42608 sw
tri 15340 42592 15348 42600 ne
rect 15348 42592 15616 42600
tri 15616 42592 15624 42600 sw
tri 15348 42584 15356 42592 ne
rect 15356 42584 15624 42592
tri 15624 42584 15632 42592 sw
tri 15356 42576 15364 42584 ne
rect 15364 42580 15632 42584
rect 15364 42576 15498 42580
tri 15364 42568 15372 42576 ne
rect 15372 42568 15498 42576
tri 15372 42560 15380 42568 ne
rect 15380 42560 15498 42568
tri 15380 42552 15388 42560 ne
rect 15388 42552 15498 42560
tri 15388 42544 15396 42552 ne
rect 15396 42544 15498 42552
tri 15396 42536 15404 42544 ne
rect 15404 42536 15498 42544
tri 15404 42528 15412 42536 ne
rect 15412 42534 15498 42536
rect 15544 42576 15632 42580
tri 15632 42576 15640 42584 sw
rect 15544 42568 15640 42576
tri 15640 42568 15648 42576 sw
rect 15544 42560 15648 42568
tri 15648 42560 15656 42568 sw
rect 15544 42552 15656 42560
tri 15656 42552 15664 42560 sw
rect 70802 42556 71000 42614
rect 15544 42544 15664 42552
tri 15664 42544 15672 42552 sw
rect 15544 42536 15672 42544
tri 15672 42536 15680 42544 sw
rect 15544 42534 15680 42536
rect 15412 42528 15680 42534
tri 15680 42528 15688 42536 sw
tri 15412 42522 15418 42528 ne
rect 15418 42527 15688 42528
tri 15688 42527 15689 42528 sw
rect 15418 42522 15689 42527
tri 15418 42514 15426 42522 ne
rect 15426 42519 15689 42522
tri 15689 42519 15697 42527 sw
rect 15426 42514 15697 42519
tri 15426 42506 15434 42514 ne
rect 15434 42511 15697 42514
tri 15697 42511 15705 42519 sw
rect 15434 42506 15705 42511
tri 15434 42498 15442 42506 ne
rect 15442 42503 15705 42506
tri 15705 42503 15713 42511 sw
rect 70802 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 15442 42498 15713 42503
tri 15442 42490 15450 42498 ne
rect 15450 42495 15713 42498
tri 15713 42495 15721 42503 sw
rect 15450 42490 15721 42495
tri 15450 42482 15458 42490 ne
rect 15458 42487 15721 42490
tri 15721 42487 15729 42495 sw
rect 15458 42482 15729 42487
tri 15458 42474 15466 42482 ne
rect 15466 42479 15729 42482
tri 15729 42479 15737 42487 sw
rect 15466 42474 15737 42479
tri 15466 42466 15474 42474 ne
rect 15474 42471 15737 42474
tri 15737 42471 15745 42479 sw
rect 15474 42466 15745 42471
tri 15474 42458 15482 42466 ne
rect 15482 42463 15745 42466
tri 15745 42463 15753 42471 sw
rect 15482 42458 15753 42463
tri 15753 42458 15758 42463 sw
tri 15482 42450 15490 42458 ne
rect 15490 42450 15758 42458
tri 15758 42450 15766 42458 sw
rect 70802 42452 71000 42510
tri 15490 42442 15498 42450 ne
rect 15498 42448 15766 42450
rect 15498 42442 15630 42448
tri 15498 42434 15506 42442 ne
rect 15506 42434 15630 42442
tri 15506 42426 15514 42434 ne
rect 15514 42426 15630 42434
tri 15514 42418 15522 42426 ne
rect 15522 42418 15630 42426
tri 15522 42410 15530 42418 ne
rect 15530 42410 15630 42418
tri 15530 42402 15538 42410 ne
rect 15538 42402 15630 42410
rect 15676 42442 15766 42448
tri 15766 42442 15774 42450 sw
rect 15676 42434 15774 42442
tri 15774 42434 15782 42442 sw
rect 15676 42426 15782 42434
tri 15782 42426 15790 42434 sw
rect 15676 42418 15790 42426
tri 15790 42418 15798 42426 sw
rect 15676 42410 15798 42418
tri 15798 42410 15806 42418 sw
rect 15676 42402 15806 42410
tri 15806 42402 15814 42410 sw
rect 70802 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
tri 15538 42401 15539 42402 ne
rect 15539 42401 15814 42402
tri 15814 42401 15815 42402 sw
tri 15539 42393 15547 42401 ne
rect 15547 42393 15815 42401
tri 15815 42393 15823 42401 sw
tri 15547 42385 15555 42393 ne
rect 15555 42385 15823 42393
tri 15823 42385 15831 42393 sw
tri 15555 42377 15563 42385 ne
rect 15563 42377 15831 42385
tri 15831 42377 15839 42385 sw
tri 15563 42369 15571 42377 ne
rect 15571 42369 15839 42377
tri 15839 42369 15847 42377 sw
tri 15571 42361 15579 42369 ne
rect 15579 42361 15847 42369
tri 15847 42361 15855 42369 sw
tri 15579 42353 15587 42361 ne
rect 15587 42353 15855 42361
tri 15855 42353 15863 42361 sw
tri 15587 42345 15595 42353 ne
rect 15595 42345 15863 42353
tri 15863 42345 15871 42353 sw
rect 70802 42348 71000 42406
tri 15595 42337 15603 42345 ne
rect 15603 42337 15871 42345
tri 15871 42337 15879 42345 sw
tri 15603 42329 15611 42337 ne
rect 15611 42329 15879 42337
tri 15879 42329 15887 42337 sw
tri 15611 42321 15619 42329 ne
rect 15619 42321 15887 42329
tri 15887 42321 15895 42329 sw
tri 15619 42313 15627 42321 ne
rect 15627 42316 15895 42321
rect 15627 42313 15762 42316
tri 15627 42305 15635 42313 ne
rect 15635 42305 15762 42313
tri 15635 42297 15643 42305 ne
rect 15643 42297 15762 42305
tri 15643 42289 15651 42297 ne
rect 15651 42289 15762 42297
tri 15651 42281 15659 42289 ne
rect 15659 42281 15762 42289
tri 15659 42273 15667 42281 ne
rect 15667 42273 15762 42281
tri 15667 42265 15675 42273 ne
rect 15675 42270 15762 42273
rect 15808 42313 15895 42316
tri 15895 42313 15903 42321 sw
rect 15808 42305 15903 42313
tri 15903 42305 15911 42313 sw
rect 15808 42297 15911 42305
tri 15911 42297 15919 42305 sw
rect 70802 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42289 15919 42297
tri 15919 42289 15927 42297 sw
rect 15808 42281 15927 42289
tri 15927 42281 15935 42289 sw
rect 15808 42273 15935 42281
tri 15935 42273 15943 42281 sw
rect 15808 42270 15943 42273
rect 15675 42265 15943 42270
tri 15943 42265 15951 42273 sw
tri 15675 42259 15681 42265 ne
rect 15681 42259 15951 42265
tri 15951 42259 15957 42265 sw
tri 15681 42251 15689 42259 ne
rect 15689 42251 15957 42259
tri 15957 42251 15965 42259 sw
tri 15689 42243 15697 42251 ne
rect 15697 42243 15965 42251
tri 15965 42243 15973 42251 sw
rect 70802 42244 71000 42302
tri 15697 42235 15705 42243 ne
rect 15705 42235 15973 42243
tri 15973 42235 15981 42243 sw
tri 15705 42227 15713 42235 ne
rect 15713 42227 15981 42235
tri 15981 42227 15989 42235 sw
tri 15713 42219 15721 42227 ne
rect 15721 42219 15989 42227
tri 15989 42219 15997 42227 sw
tri 15721 42211 15729 42219 ne
rect 15729 42211 15997 42219
tri 15997 42211 16005 42219 sw
tri 15729 42203 15737 42211 ne
rect 15737 42203 16005 42211
tri 16005 42203 16013 42211 sw
tri 15737 42195 15745 42203 ne
rect 15745 42195 16013 42203
tri 16013 42195 16021 42203 sw
rect 70802 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
tri 15745 42187 15753 42195 ne
rect 15753 42187 16021 42195
tri 16021 42187 16029 42195 sw
tri 15753 42179 15761 42187 ne
rect 15761 42184 16029 42187
rect 15761 42179 15894 42184
tri 15761 42171 15769 42179 ne
rect 15769 42171 15894 42179
tri 15769 42163 15777 42171 ne
rect 15777 42163 15894 42171
tri 15777 42155 15785 42163 ne
rect 15785 42155 15894 42163
tri 15785 42147 15793 42155 ne
rect 15793 42147 15894 42155
tri 15793 42139 15801 42147 ne
rect 15801 42139 15894 42147
tri 15801 42131 15809 42139 ne
rect 15809 42138 15894 42139
rect 15940 42179 16029 42184
tri 16029 42179 16037 42187 sw
rect 15940 42171 16037 42179
tri 16037 42171 16045 42179 sw
rect 15940 42163 16045 42171
tri 16045 42163 16053 42171 sw
rect 15940 42155 16053 42163
tri 16053 42155 16061 42163 sw
rect 15940 42147 16061 42155
tri 16061 42147 16069 42155 sw
rect 15940 42139 16069 42147
tri 16069 42139 16077 42147 sw
rect 70802 42140 71000 42198
rect 15940 42138 16077 42139
rect 15809 42131 16077 42138
tri 16077 42131 16085 42139 sw
tri 15809 42125 15815 42131 ne
rect 15815 42125 16085 42131
tri 16085 42125 16091 42131 sw
tri 15815 42117 15823 42125 ne
rect 15823 42117 16091 42125
tri 16091 42117 16099 42125 sw
tri 15823 42109 15831 42117 ne
rect 15831 42109 16099 42117
tri 16099 42109 16107 42117 sw
tri 15831 42101 15839 42109 ne
rect 15839 42101 16107 42109
tri 16107 42101 16115 42109 sw
tri 15839 42093 15847 42101 ne
rect 15847 42093 16115 42101
tri 16115 42093 16123 42101 sw
rect 70802 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15847 42085 15855 42093 ne
rect 15855 42085 16123 42093
tri 16123 42085 16131 42093 sw
tri 15855 42077 15863 42085 ne
rect 15863 42077 16131 42085
tri 16131 42077 16139 42085 sw
tri 15863 42069 15871 42077 ne
rect 15871 42069 16139 42077
tri 16139 42069 16147 42077 sw
tri 15871 42061 15879 42069 ne
rect 15879 42061 16147 42069
tri 16147 42061 16155 42069 sw
tri 15879 42053 15887 42061 ne
rect 15887 42053 16155 42061
tri 16155 42053 16163 42061 sw
tri 15887 42045 15895 42053 ne
rect 15895 42052 16163 42053
rect 15895 42045 16026 42052
tri 15895 42037 15903 42045 ne
rect 15903 42037 16026 42045
tri 15903 42029 15911 42037 ne
rect 15911 42029 16026 42037
tri 15911 42021 15919 42029 ne
rect 15919 42021 16026 42029
tri 15919 42013 15927 42021 ne
rect 15927 42013 16026 42021
tri 15927 42005 15935 42013 ne
rect 15935 42006 16026 42013
rect 16072 42045 16163 42052
tri 16163 42045 16171 42053 sw
rect 16072 42037 16171 42045
tri 16171 42037 16179 42045 sw
rect 16072 42029 16179 42037
tri 16179 42029 16187 42037 sw
rect 70802 42036 71000 42094
rect 16072 42021 16187 42029
tri 16187 42021 16195 42029 sw
rect 16072 42013 16195 42021
tri 16195 42013 16203 42021 sw
rect 16072 42010 16203 42013
tri 16203 42010 16206 42013 sw
rect 16072 42006 16206 42010
rect 15935 42005 16206 42006
tri 15935 42002 15938 42005 ne
rect 15938 42002 16206 42005
tri 16206 42002 16214 42010 sw
tri 15938 41994 15946 42002 ne
rect 15946 41994 16214 42002
tri 16214 41994 16222 42002 sw
tri 15946 41986 15954 41994 ne
rect 15954 41986 16222 41994
tri 16222 41986 16230 41994 sw
rect 70802 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15954 41978 15962 41986 ne
rect 15962 41978 16230 41986
tri 16230 41978 16238 41986 sw
tri 15962 41970 15970 41978 ne
rect 15970 41970 16238 41978
tri 16238 41970 16246 41978 sw
tri 15970 41962 15978 41970 ne
rect 15978 41962 16246 41970
tri 16246 41962 16254 41970 sw
tri 15978 41954 15986 41962 ne
rect 15986 41954 16254 41962
tri 16254 41954 16262 41962 sw
tri 15986 41946 15994 41954 ne
rect 15994 41946 16262 41954
tri 16262 41946 16270 41954 sw
tri 15994 41938 16002 41946 ne
rect 16002 41938 16270 41946
tri 16270 41938 16278 41946 sw
tri 16002 41930 16010 41938 ne
rect 16010 41930 16278 41938
tri 16278 41930 16286 41938 sw
rect 70802 41932 71000 41990
tri 16010 41922 16018 41930 ne
rect 16018 41922 16286 41930
tri 16286 41922 16294 41930 sw
tri 16018 41914 16026 41922 ne
rect 16026 41920 16294 41922
rect 16026 41914 16158 41920
tri 16026 41906 16034 41914 ne
rect 16034 41906 16158 41914
tri 16034 41898 16042 41906 ne
rect 16042 41898 16158 41906
tri 16042 41890 16050 41898 ne
rect 16050 41890 16158 41898
tri 16050 41882 16058 41890 ne
rect 16058 41882 16158 41890
tri 16058 41874 16066 41882 ne
rect 16066 41874 16158 41882
rect 16204 41914 16294 41920
tri 16294 41914 16302 41922 sw
rect 16204 41906 16302 41914
tri 16302 41906 16310 41914 sw
rect 16204 41898 16310 41906
tri 16310 41898 16318 41906 sw
rect 16204 41890 16318 41898
tri 16318 41890 16326 41898 sw
rect 16204 41882 16326 41890
tri 16326 41882 16334 41890 sw
rect 70802 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 16204 41874 16334 41882
tri 16334 41874 16342 41882 sw
tri 16066 41866 16074 41874 ne
rect 16074 41866 16342 41874
tri 16342 41866 16350 41874 sw
tri 16074 41865 16075 41866 ne
rect 16075 41865 16350 41866
tri 16350 41865 16351 41866 sw
tri 16075 41857 16083 41865 ne
rect 16083 41857 16351 41865
tri 16351 41857 16359 41865 sw
tri 16083 41849 16091 41857 ne
rect 16091 41849 16359 41857
tri 16359 41849 16367 41857 sw
tri 16091 41841 16099 41849 ne
rect 16099 41841 16367 41849
tri 16367 41841 16375 41849 sw
tri 16099 41833 16107 41841 ne
rect 16107 41833 16375 41841
tri 16375 41833 16383 41841 sw
tri 16107 41825 16115 41833 ne
rect 16115 41825 16383 41833
tri 16383 41825 16391 41833 sw
rect 70802 41828 71000 41886
tri 16115 41817 16123 41825 ne
rect 16123 41817 16391 41825
tri 16391 41817 16399 41825 sw
tri 16123 41809 16131 41817 ne
rect 16131 41809 16399 41817
tri 16399 41809 16407 41817 sw
tri 16131 41801 16139 41809 ne
rect 16139 41801 16407 41809
tri 16407 41801 16415 41809 sw
tri 16139 41793 16147 41801 ne
rect 16147 41793 16415 41801
tri 16415 41793 16423 41801 sw
tri 16147 41785 16155 41793 ne
rect 16155 41788 16423 41793
rect 16155 41785 16290 41788
tri 16155 41777 16163 41785 ne
rect 16163 41777 16290 41785
tri 16163 41769 16171 41777 ne
rect 16171 41769 16290 41777
tri 16171 41761 16179 41769 ne
rect 16179 41761 16290 41769
tri 16179 41753 16187 41761 ne
rect 16187 41753 16290 41761
tri 16187 41745 16195 41753 ne
rect 16195 41745 16290 41753
tri 16195 41737 16203 41745 ne
rect 16203 41742 16290 41745
rect 16336 41785 16423 41788
tri 16423 41785 16431 41793 sw
rect 16336 41777 16431 41785
tri 16431 41777 16439 41785 sw
rect 70802 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41769 16439 41777
tri 16439 41769 16447 41777 sw
rect 16336 41761 16447 41769
tri 16447 41761 16455 41769 sw
rect 16336 41753 16455 41761
tri 16455 41753 16463 41761 sw
rect 16336 41745 16463 41753
tri 16463 41745 16471 41753 sw
rect 16336 41742 16471 41745
rect 16203 41737 16471 41742
tri 16471 41737 16479 41745 sw
tri 16203 41729 16211 41737 ne
rect 16211 41731 16479 41737
tri 16479 41731 16485 41737 sw
rect 16211 41729 16485 41731
tri 16211 41726 16214 41729 ne
rect 16214 41726 16485 41729
tri 16214 41718 16222 41726 ne
rect 16222 41723 16485 41726
tri 16485 41723 16493 41731 sw
rect 70802 41724 71000 41782
rect 16222 41718 16493 41723
tri 16222 41710 16230 41718 ne
rect 16230 41715 16493 41718
tri 16493 41715 16501 41723 sw
rect 16230 41710 16501 41715
tri 16230 41702 16238 41710 ne
rect 16238 41707 16501 41710
tri 16501 41707 16509 41715 sw
rect 16238 41702 16509 41707
tri 16238 41694 16246 41702 ne
rect 16246 41699 16509 41702
tri 16509 41699 16517 41707 sw
rect 16246 41694 16517 41699
tri 16246 41686 16254 41694 ne
rect 16254 41691 16517 41694
tri 16517 41691 16525 41699 sw
rect 16254 41686 16525 41691
tri 16254 41678 16262 41686 ne
rect 16262 41683 16525 41686
tri 16525 41683 16533 41691 sw
rect 16262 41678 16533 41683
tri 16262 41670 16270 41678 ne
rect 16270 41675 16533 41678
tri 16533 41675 16541 41683 sw
rect 70802 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16270 41670 16541 41675
tri 16270 41662 16278 41670 ne
rect 16278 41667 16541 41670
tri 16541 41667 16549 41675 sw
rect 16278 41662 16549 41667
tri 16278 41654 16286 41662 ne
rect 16286 41659 16549 41662
tri 16549 41659 16557 41667 sw
rect 16286 41656 16557 41659
rect 16286 41654 16422 41656
tri 16286 41646 16294 41654 ne
rect 16294 41646 16422 41654
tri 16294 41638 16302 41646 ne
rect 16302 41638 16422 41646
tri 16302 41630 16310 41638 ne
rect 16310 41630 16422 41638
tri 16310 41622 16318 41630 ne
rect 16318 41622 16422 41630
tri 16318 41614 16326 41622 ne
rect 16326 41614 16422 41622
tri 16326 41606 16334 41614 ne
rect 16334 41610 16422 41614
rect 16468 41651 16557 41656
tri 16557 41651 16565 41659 sw
rect 16468 41643 16565 41651
tri 16565 41643 16573 41651 sw
rect 16468 41635 16573 41643
tri 16573 41635 16581 41643 sw
rect 16468 41627 16581 41635
tri 16581 41627 16589 41635 sw
rect 16468 41619 16589 41627
tri 16589 41619 16597 41627 sw
rect 70802 41620 71000 41678
rect 16468 41611 16597 41619
tri 16597 41611 16605 41619 sw
rect 16468 41610 16605 41611
rect 16334 41606 16605 41610
tri 16334 41598 16342 41606 ne
rect 16342 41603 16605 41606
tri 16605 41603 16613 41611 sw
rect 16342 41598 16613 41603
tri 16342 41590 16350 41598 ne
rect 16350 41595 16613 41598
tri 16613 41595 16621 41603 sw
rect 16350 41590 16621 41595
tri 16350 41589 16351 41590 ne
rect 16351 41589 16621 41590
tri 16621 41589 16627 41595 sw
tri 16351 41581 16359 41589 ne
rect 16359 41581 16627 41589
tri 16627 41581 16635 41589 sw
tri 16359 41573 16367 41581 ne
rect 16367 41573 16635 41581
tri 16635 41573 16643 41581 sw
rect 70802 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16367 41565 16375 41573 ne
rect 16375 41565 16643 41573
tri 16643 41565 16651 41573 sw
tri 16375 41557 16383 41565 ne
rect 16383 41557 16651 41565
tri 16651 41557 16659 41565 sw
tri 16383 41549 16391 41557 ne
rect 16391 41549 16659 41557
tri 16659 41549 16667 41557 sw
tri 16391 41541 16399 41549 ne
rect 16399 41541 16667 41549
tri 16667 41541 16675 41549 sw
tri 16399 41533 16407 41541 ne
rect 16407 41533 16675 41541
tri 16675 41533 16683 41541 sw
tri 16407 41525 16415 41533 ne
rect 16415 41525 16683 41533
tri 16683 41525 16691 41533 sw
tri 16415 41517 16423 41525 ne
rect 16423 41524 16691 41525
rect 16423 41517 16554 41524
tri 16423 41509 16431 41517 ne
rect 16431 41509 16554 41517
tri 16431 41501 16439 41509 ne
rect 16439 41501 16554 41509
tri 16439 41493 16447 41501 ne
rect 16447 41493 16554 41501
tri 16447 41485 16455 41493 ne
rect 16455 41485 16554 41493
tri 16455 41477 16463 41485 ne
rect 16463 41478 16554 41485
rect 16600 41517 16691 41524
tri 16691 41517 16699 41525 sw
rect 16600 41509 16699 41517
tri 16699 41509 16707 41517 sw
rect 70802 41516 71000 41574
rect 16600 41501 16707 41509
tri 16707 41501 16715 41509 sw
rect 16600 41493 16715 41501
tri 16715 41493 16723 41501 sw
rect 16600 41485 16723 41493
tri 16723 41485 16731 41493 sw
rect 16600 41479 16731 41485
tri 16731 41479 16737 41485 sw
rect 16600 41478 16737 41479
rect 16463 41477 16737 41478
tri 16463 41469 16471 41477 ne
rect 16471 41471 16737 41477
tri 16737 41471 16745 41479 sw
rect 16471 41469 16745 41471
tri 16471 41465 16475 41469 ne
rect 16475 41465 16745 41469
tri 16475 41457 16483 41465 ne
rect 16483 41463 16745 41465
tri 16745 41463 16753 41471 sw
rect 70802 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 16483 41457 16753 41463
tri 16483 41449 16491 41457 ne
rect 16491 41455 16753 41457
tri 16753 41455 16761 41463 sw
rect 16491 41449 16761 41455
tri 16491 41441 16499 41449 ne
rect 16499 41447 16761 41449
tri 16761 41447 16769 41455 sw
rect 16499 41441 16769 41447
tri 16499 41433 16507 41441 ne
rect 16507 41439 16769 41441
tri 16769 41439 16777 41447 sw
rect 16507 41433 16777 41439
tri 16507 41425 16515 41433 ne
rect 16515 41431 16777 41433
tri 16777 41431 16785 41439 sw
rect 16515 41425 16785 41431
tri 16515 41417 16523 41425 ne
rect 16523 41423 16785 41425
tri 16785 41423 16793 41431 sw
rect 16523 41417 16793 41423
tri 16523 41409 16531 41417 ne
rect 16531 41415 16793 41417
tri 16793 41415 16801 41423 sw
rect 16531 41409 16801 41415
tri 16531 41401 16539 41409 ne
rect 16539 41407 16801 41409
tri 16801 41407 16809 41415 sw
rect 70802 41412 71000 41470
rect 16539 41401 16809 41407
tri 16539 41393 16547 41401 ne
rect 16547 41399 16809 41401
tri 16809 41399 16817 41407 sw
rect 16547 41393 16817 41399
tri 16547 41385 16555 41393 ne
rect 16555 41392 16817 41393
rect 16555 41385 16686 41392
tri 16555 41377 16563 41385 ne
rect 16563 41377 16686 41385
tri 16563 41369 16571 41377 ne
rect 16571 41369 16686 41377
tri 16571 41361 16579 41369 ne
rect 16579 41361 16686 41369
tri 16579 41353 16587 41361 ne
rect 16587 41353 16686 41361
tri 16587 41345 16595 41353 ne
rect 16595 41346 16686 41353
rect 16732 41391 16817 41392
tri 16817 41391 16825 41399 sw
rect 16732 41383 16825 41391
tri 16825 41383 16833 41391 sw
rect 16732 41375 16833 41383
tri 16833 41375 16841 41383 sw
rect 16732 41367 16841 41375
tri 16841 41367 16849 41375 sw
rect 16732 41359 16849 41367
tri 16849 41359 16857 41367 sw
rect 70802 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 16732 41358 16857 41359
tri 16857 41358 16858 41359 sw
rect 16732 41350 16858 41358
tri 16858 41350 16866 41358 sw
rect 16732 41346 16866 41350
rect 16595 41345 16866 41346
tri 16595 41337 16603 41345 ne
rect 16603 41342 16866 41345
tri 16866 41342 16874 41350 sw
rect 16603 41337 16874 41342
tri 16603 41329 16611 41337 ne
rect 16611 41334 16874 41337
tri 16874 41334 16882 41342 sw
rect 16611 41329 16882 41334
tri 16611 41326 16614 41329 ne
rect 16614 41326 16882 41329
tri 16882 41326 16890 41334 sw
tri 16614 41318 16622 41326 ne
rect 16622 41318 16890 41326
tri 16890 41318 16898 41326 sw
tri 16622 41310 16630 41318 ne
rect 16630 41310 16898 41318
tri 16898 41310 16906 41318 sw
tri 16630 41302 16638 41310 ne
rect 16638 41302 16906 41310
tri 16906 41302 16914 41310 sw
rect 70802 41308 71000 41366
tri 16638 41294 16646 41302 ne
rect 16646 41294 16914 41302
tri 16914 41294 16922 41302 sw
tri 16646 41286 16654 41294 ne
rect 16654 41286 16922 41294
tri 16922 41286 16930 41294 sw
tri 16654 41278 16662 41286 ne
rect 16662 41278 16930 41286
tri 16930 41278 16938 41286 sw
tri 16662 41270 16670 41278 ne
rect 16670 41270 16938 41278
tri 16938 41270 16946 41278 sw
tri 16670 41262 16678 41270 ne
rect 16678 41262 16946 41270
tri 16946 41262 16954 41270 sw
rect 70802 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
tri 16678 41254 16686 41262 ne
rect 16686 41260 16954 41262
rect 16686 41254 16818 41260
tri 16686 41246 16694 41254 ne
rect 16694 41246 16818 41254
tri 16694 41239 16701 41246 ne
rect 16701 41239 16818 41246
tri 16701 41231 16709 41239 ne
rect 16709 41231 16818 41239
tri 16709 41223 16717 41231 ne
rect 16717 41223 16818 41231
tri 16717 41215 16725 41223 ne
rect 16725 41215 16818 41223
tri 16725 41207 16733 41215 ne
rect 16733 41214 16818 41215
rect 16864 41255 16954 41260
tri 16954 41255 16961 41262 sw
rect 16864 41247 16961 41255
tri 16961 41247 16969 41255 sw
rect 16864 41239 16969 41247
tri 16969 41239 16977 41247 sw
rect 16864 41231 16977 41239
tri 16977 41231 16985 41239 sw
rect 16864 41223 16985 41231
tri 16985 41223 16993 41231 sw
rect 16864 41215 16993 41223
tri 16993 41215 17001 41223 sw
rect 16864 41214 17001 41215
rect 16733 41207 17001 41214
tri 17001 41207 17009 41215 sw
tri 16733 41199 16741 41207 ne
rect 16741 41199 17009 41207
tri 17009 41199 17017 41207 sw
rect 70802 41204 71000 41262
tri 16741 41191 16749 41199 ne
rect 16749 41191 17017 41199
tri 17017 41191 17025 41199 sw
tri 16749 41183 16757 41191 ne
rect 16757 41189 17025 41191
tri 17025 41189 17027 41191 sw
rect 16757 41183 17027 41189
tri 16757 41178 16762 41183 ne
rect 16762 41181 17027 41183
tri 17027 41181 17035 41189 sw
rect 16762 41178 17035 41181
tri 16762 41170 16770 41178 ne
rect 16770 41173 17035 41178
tri 17035 41173 17043 41181 sw
rect 16770 41170 17043 41173
tri 16770 41162 16778 41170 ne
rect 16778 41165 17043 41170
tri 17043 41165 17051 41173 sw
rect 16778 41162 17051 41165
tri 16778 41154 16786 41162 ne
rect 16786 41157 17051 41162
tri 17051 41157 17059 41165 sw
rect 70802 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
rect 16786 41154 17059 41157
tri 16786 41146 16794 41154 ne
rect 16794 41149 17059 41154
tri 17059 41149 17067 41157 sw
rect 16794 41146 17067 41149
tri 16794 41138 16802 41146 ne
rect 16802 41141 17067 41146
tri 17067 41141 17075 41149 sw
rect 16802 41138 17075 41141
tri 16802 41130 16810 41138 ne
rect 16810 41133 17075 41138
tri 17075 41133 17083 41141 sw
rect 16810 41130 17083 41133
tri 16810 41122 16818 41130 ne
rect 16818 41128 17083 41130
rect 16818 41122 16950 41128
tri 16818 41114 16826 41122 ne
rect 16826 41114 16950 41122
tri 16826 41106 16834 41114 ne
rect 16834 41106 16950 41114
tri 16834 41098 16842 41106 ne
rect 16842 41098 16950 41106
tri 16842 41090 16850 41098 ne
rect 16850 41090 16950 41098
tri 16850 41082 16858 41090 ne
rect 16858 41082 16950 41090
rect 16996 41125 17083 41128
tri 17083 41125 17091 41133 sw
rect 16996 41117 17091 41125
tri 17091 41117 17099 41125 sw
rect 16996 41109 17099 41117
tri 17099 41109 17107 41117 sw
rect 16996 41101 17107 41109
tri 17107 41101 17115 41109 sw
rect 16996 41093 17115 41101
tri 17115 41093 17123 41101 sw
rect 70802 41100 71000 41158
rect 16996 41085 17123 41093
tri 17123 41085 17131 41093 sw
rect 16996 41082 17131 41085
tri 16858 41074 16866 41082 ne
rect 16866 41077 17131 41082
tri 17131 41077 17139 41085 sw
rect 16866 41074 17139 41077
tri 16866 41066 16874 41074 ne
rect 16874 41069 17139 41074
tri 17139 41069 17147 41077 sw
rect 16874 41066 17147 41069
tri 16874 41058 16882 41066 ne
rect 16882 41061 17147 41066
tri 17147 41061 17155 41069 sw
rect 16882 41058 17155 41061
tri 16882 41050 16890 41058 ne
rect 16890 41053 17155 41058
tri 17155 41053 17163 41061 sw
rect 70802 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 16890 41050 17163 41053
tri 16890 41042 16898 41050 ne
rect 16898 41045 17163 41050
tri 17163 41045 17171 41053 sw
rect 16898 41043 17171 41045
tri 17171 41043 17173 41045 sw
rect 16898 41042 17173 41043
tri 16898 41035 16905 41042 ne
rect 16905 41035 17173 41042
tri 17173 41035 17181 41043 sw
tri 16905 41027 16913 41035 ne
rect 16913 41027 17181 41035
tri 17181 41027 17189 41035 sw
tri 16913 41019 16921 41027 ne
rect 16921 41019 17189 41027
tri 17189 41019 17197 41027 sw
tri 16921 41011 16929 41019 ne
rect 16929 41011 17197 41019
tri 17197 41011 17205 41019 sw
tri 16929 41003 16937 41011 ne
rect 16937 41003 17205 41011
tri 17205 41003 17213 41011 sw
tri 16937 40995 16945 41003 ne
rect 16945 40996 17213 41003
rect 16945 40995 17082 40996
tri 16945 40987 16953 40995 ne
rect 16953 40987 17082 40995
tri 16953 40979 16961 40987 ne
rect 16961 40979 17082 40987
tri 16961 40971 16969 40979 ne
rect 16969 40971 17082 40979
tri 16969 40963 16977 40971 ne
rect 16977 40963 17082 40971
tri 16977 40955 16985 40963 ne
rect 16985 40955 17082 40963
tri 16985 40947 16993 40955 ne
rect 16993 40950 17082 40955
rect 17128 40995 17213 40996
tri 17213 40995 17221 41003 sw
rect 70802 40996 71000 41054
rect 17128 40987 17221 40995
tri 17221 40987 17229 40995 sw
rect 17128 40979 17229 40987
tri 17229 40979 17237 40987 sw
rect 17128 40971 17237 40979
tri 17237 40971 17245 40979 sw
rect 17128 40963 17245 40971
tri 17245 40963 17253 40971 sw
rect 17128 40955 17253 40963
tri 17253 40955 17261 40963 sw
rect 17128 40950 17261 40955
rect 16993 40947 17261 40950
tri 17261 40947 17269 40955 sw
rect 70802 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
tri 16993 40939 17001 40947 ne
rect 17001 40939 17269 40947
tri 17269 40939 17277 40947 sw
tri 17001 40931 17009 40939 ne
rect 17009 40931 17277 40939
tri 17277 40931 17285 40939 sw
tri 17009 40923 17017 40931 ne
rect 17017 40923 17285 40931
tri 17285 40923 17293 40931 sw
tri 17017 40915 17025 40923 ne
rect 17025 40915 17293 40923
tri 17293 40915 17301 40923 sw
tri 17025 40907 17033 40915 ne
rect 17033 40907 17301 40915
tri 17301 40907 17309 40915 sw
tri 17033 40905 17035 40907 ne
rect 17035 40905 17309 40907
tri 17309 40905 17311 40907 sw
tri 17035 40897 17043 40905 ne
rect 17043 40897 17311 40905
tri 17311 40897 17319 40905 sw
tri 17043 40889 17051 40897 ne
rect 17051 40889 17319 40897
tri 17319 40889 17327 40897 sw
rect 70802 40892 71000 40950
tri 17051 40881 17059 40889 ne
rect 17059 40881 17327 40889
tri 17327 40881 17335 40889 sw
tri 17059 40873 17067 40881 ne
rect 17067 40873 17335 40881
tri 17335 40873 17343 40881 sw
tri 17067 40865 17075 40873 ne
rect 17075 40865 17343 40873
tri 17343 40865 17351 40873 sw
tri 17075 40857 17083 40865 ne
rect 17083 40864 17351 40865
rect 17083 40857 17214 40864
tri 17083 40849 17091 40857 ne
rect 17091 40849 17214 40857
tri 17091 40841 17099 40849 ne
rect 17099 40841 17214 40849
tri 17099 40833 17107 40841 ne
rect 17107 40833 17214 40841
tri 17107 40825 17115 40833 ne
rect 17115 40825 17214 40833
tri 17115 40817 17123 40825 ne
rect 17123 40818 17214 40825
rect 17260 40857 17351 40864
tri 17351 40857 17359 40865 sw
rect 17260 40849 17359 40857
tri 17359 40849 17367 40857 sw
rect 17260 40841 17367 40849
tri 17367 40841 17375 40849 sw
rect 70802 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40833 17375 40841
tri 17375 40833 17383 40841 sw
rect 17260 40825 17383 40833
tri 17383 40825 17391 40833 sw
rect 17260 40818 17391 40825
rect 17123 40817 17391 40818
tri 17391 40817 17399 40825 sw
tri 17123 40809 17131 40817 ne
rect 17131 40814 17399 40817
tri 17399 40814 17402 40817 sw
rect 17131 40809 17402 40814
tri 17131 40801 17139 40809 ne
rect 17139 40806 17402 40809
tri 17402 40806 17410 40814 sw
rect 17139 40801 17410 40806
tri 17139 40793 17147 40801 ne
rect 17147 40798 17410 40801
tri 17410 40798 17418 40806 sw
rect 17147 40793 17418 40798
tri 17147 40785 17155 40793 ne
rect 17155 40790 17418 40793
tri 17418 40790 17426 40798 sw
rect 17155 40785 17426 40790
tri 17155 40777 17163 40785 ne
rect 17163 40782 17426 40785
tri 17426 40782 17434 40790 sw
rect 70802 40788 71000 40846
rect 17163 40777 17434 40782
tri 17163 40771 17169 40777 ne
rect 17169 40774 17434 40777
tri 17434 40774 17442 40782 sw
rect 17169 40771 17442 40774
tri 17169 40763 17177 40771 ne
rect 17177 40766 17442 40771
tri 17442 40766 17450 40774 sw
rect 17177 40763 17450 40766
tri 17177 40755 17185 40763 ne
rect 17185 40758 17450 40763
tri 17450 40758 17458 40766 sw
rect 17185 40755 17458 40758
tri 17185 40747 17193 40755 ne
rect 17193 40750 17458 40755
tri 17458 40750 17466 40758 sw
rect 17193 40747 17466 40750
tri 17193 40739 17201 40747 ne
rect 17201 40742 17466 40747
tri 17466 40742 17474 40750 sw
rect 70802 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17201 40739 17474 40742
tri 17201 40731 17209 40739 ne
rect 17209 40734 17474 40739
tri 17474 40734 17482 40742 sw
rect 17209 40732 17482 40734
rect 17209 40731 17346 40732
tri 17209 40723 17217 40731 ne
rect 17217 40723 17346 40731
tri 17217 40715 17225 40723 ne
rect 17225 40715 17346 40723
tri 17225 40707 17233 40715 ne
rect 17233 40707 17346 40715
tri 17233 40699 17241 40707 ne
rect 17241 40699 17346 40707
tri 17241 40691 17249 40699 ne
rect 17249 40691 17346 40699
tri 17249 40683 17257 40691 ne
rect 17257 40686 17346 40691
rect 17392 40726 17482 40732
tri 17482 40726 17490 40734 sw
rect 17392 40719 17490 40726
tri 17490 40719 17497 40726 sw
rect 17392 40711 17497 40719
tri 17497 40711 17505 40719 sw
rect 17392 40703 17505 40711
tri 17505 40703 17513 40711 sw
rect 17392 40695 17513 40703
tri 17513 40695 17521 40703 sw
rect 17392 40687 17521 40695
tri 17521 40687 17529 40695 sw
rect 17392 40686 17529 40687
rect 17257 40683 17529 40686
tri 17529 40683 17533 40687 sw
rect 70802 40684 71000 40742
tri 17257 40675 17265 40683 ne
rect 17265 40675 17533 40683
tri 17533 40675 17541 40683 sw
tri 17265 40667 17273 40675 ne
rect 17273 40667 17541 40675
tri 17541 40667 17549 40675 sw
tri 17273 40659 17281 40667 ne
rect 17281 40659 17549 40667
tri 17549 40659 17557 40667 sw
tri 17281 40651 17289 40659 ne
rect 17289 40651 17557 40659
tri 17557 40651 17565 40659 sw
tri 17289 40643 17297 40651 ne
rect 17297 40643 17565 40651
tri 17565 40643 17573 40651 sw
tri 17297 40635 17305 40643 ne
rect 17305 40635 17573 40643
tri 17573 40635 17581 40643 sw
rect 70802 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17305 40631 17309 40635 ne
rect 17309 40631 17581 40635
tri 17309 40623 17317 40631 ne
rect 17317 40627 17581 40631
tri 17581 40627 17589 40635 sw
rect 17317 40623 17589 40627
tri 17317 40615 17325 40623 ne
rect 17325 40619 17589 40623
tri 17589 40619 17597 40627 sw
rect 17325 40615 17597 40619
tri 17325 40607 17333 40615 ne
rect 17333 40611 17597 40615
tri 17597 40611 17605 40619 sw
rect 17333 40607 17605 40611
tri 17333 40599 17341 40607 ne
rect 17341 40603 17605 40607
tri 17605 40603 17613 40611 sw
rect 17341 40600 17613 40603
rect 17341 40599 17478 40600
tri 17341 40591 17349 40599 ne
rect 17349 40591 17478 40599
tri 17349 40583 17357 40591 ne
rect 17357 40583 17478 40591
tri 17357 40575 17365 40583 ne
rect 17365 40575 17478 40583
tri 17365 40567 17373 40575 ne
rect 17373 40567 17478 40575
tri 17373 40559 17381 40567 ne
rect 17381 40559 17478 40567
tri 17381 40551 17389 40559 ne
rect 17389 40554 17478 40559
rect 17524 40595 17613 40600
tri 17613 40595 17621 40603 sw
rect 17524 40587 17621 40595
tri 17621 40587 17629 40595 sw
rect 17524 40579 17629 40587
tri 17629 40579 17637 40587 sw
rect 70802 40580 71000 40638
rect 17524 40571 17637 40579
tri 17637 40571 17645 40579 sw
rect 17524 40566 17645 40571
tri 17645 40566 17650 40571 sw
rect 17524 40558 17650 40566
tri 17650 40558 17658 40566 sw
rect 17524 40554 17658 40558
rect 17389 40551 17658 40554
tri 17389 40543 17397 40551 ne
rect 17397 40550 17658 40551
tri 17658 40550 17666 40558 sw
rect 17397 40543 17666 40550
tri 17397 40535 17405 40543 ne
rect 17405 40542 17666 40543
tri 17666 40542 17674 40550 sw
rect 17405 40535 17674 40542
tri 17405 40534 17406 40535 ne
rect 17406 40534 17674 40535
tri 17674 40534 17682 40542 sw
rect 70802 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17406 40526 17414 40534 ne
rect 17414 40526 17682 40534
tri 17682 40526 17690 40534 sw
tri 17414 40518 17422 40526 ne
rect 17422 40518 17690 40526
tri 17690 40518 17698 40526 sw
tri 17422 40510 17430 40518 ne
rect 17430 40510 17698 40518
tri 17698 40510 17706 40518 sw
tri 17430 40502 17438 40510 ne
rect 17438 40502 17706 40510
tri 17706 40502 17714 40510 sw
tri 17438 40494 17446 40502 ne
rect 17446 40494 17714 40502
tri 17714 40494 17722 40502 sw
tri 17446 40486 17454 40494 ne
rect 17454 40486 17722 40494
tri 17722 40486 17730 40494 sw
tri 17454 40478 17462 40486 ne
rect 17462 40478 17730 40486
tri 17730 40478 17738 40486 sw
tri 17462 40470 17470 40478 ne
rect 17470 40470 17738 40478
tri 17738 40470 17746 40478 sw
rect 70802 40476 71000 40534
tri 17470 40462 17478 40470 ne
rect 17478 40468 17746 40470
rect 17478 40462 17610 40468
tri 17478 40454 17486 40462 ne
rect 17486 40454 17610 40462
tri 17486 40446 17494 40454 ne
rect 17494 40446 17610 40454
tri 17494 40443 17497 40446 ne
rect 17497 40443 17610 40446
tri 17497 40435 17505 40443 ne
rect 17505 40435 17610 40443
tri 17505 40427 17513 40435 ne
rect 17513 40427 17610 40435
tri 17513 40419 17521 40427 ne
rect 17521 40422 17610 40427
rect 17656 40462 17746 40468
tri 17746 40462 17754 40470 sw
rect 17656 40454 17754 40462
tri 17754 40454 17762 40462 sw
rect 17656 40446 17762 40454
tri 17762 40446 17770 40454 sw
rect 17656 40443 17770 40446
tri 17770 40443 17773 40446 sw
rect 17656 40435 17773 40443
tri 17773 40435 17781 40443 sw
rect 17656 40427 17781 40435
tri 17781 40427 17789 40435 sw
rect 70802 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 17656 40422 17789 40427
rect 17521 40419 17789 40422
tri 17789 40419 17797 40427 sw
tri 17521 40411 17529 40419 ne
rect 17529 40411 17797 40419
tri 17797 40411 17805 40419 sw
tri 17529 40403 17537 40411 ne
rect 17537 40403 17805 40411
tri 17805 40403 17813 40411 sw
tri 17537 40395 17545 40403 ne
rect 17545 40395 17813 40403
tri 17813 40395 17821 40403 sw
tri 17545 40387 17553 40395 ne
rect 17553 40387 17821 40395
tri 17821 40387 17829 40395 sw
tri 17553 40379 17561 40387 ne
rect 17561 40379 17829 40387
tri 17829 40379 17837 40387 sw
tri 17561 40371 17569 40379 ne
rect 17569 40371 17837 40379
tri 17837 40371 17845 40379 sw
rect 70802 40372 71000 40430
tri 17569 40363 17577 40371 ne
rect 17577 40363 17845 40371
tri 17845 40363 17853 40371 sw
tri 17577 40355 17585 40363 ne
rect 17585 40355 17853 40363
tri 17853 40355 17861 40363 sw
tri 17585 40347 17593 40355 ne
rect 17593 40347 17861 40355
tri 17861 40347 17869 40355 sw
tri 17593 40339 17601 40347 ne
rect 17601 40339 17869 40347
tri 17869 40339 17877 40347 sw
tri 17601 40331 17609 40339 ne
rect 17609 40336 17877 40339
rect 17609 40331 17742 40336
tri 17609 40323 17617 40331 ne
rect 17617 40323 17742 40331
tri 17617 40316 17624 40323 ne
rect 17624 40316 17742 40323
tri 17624 40308 17632 40316 ne
rect 17632 40308 17742 40316
tri 17632 40300 17640 40308 ne
rect 17640 40300 17742 40308
tri 17640 40292 17648 40300 ne
rect 17648 40292 17742 40300
tri 17648 40284 17656 40292 ne
rect 17656 40290 17742 40292
rect 17788 40331 17877 40336
tri 17877 40331 17885 40339 sw
rect 17788 40323 17885 40331
tri 17885 40323 17893 40331 sw
rect 70802 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17788 40319 17893 40323
tri 17893 40319 17897 40323 sw
rect 17788 40311 17897 40319
tri 17897 40311 17905 40319 sw
rect 17788 40303 17905 40311
tri 17905 40303 17913 40311 sw
rect 17788 40295 17913 40303
tri 17913 40295 17921 40303 sw
rect 17788 40290 17921 40295
rect 17656 40287 17921 40290
tri 17921 40287 17929 40295 sw
rect 17656 40284 17929 40287
tri 17656 40276 17664 40284 ne
rect 17664 40279 17929 40284
tri 17929 40279 17937 40287 sw
rect 17664 40276 17937 40279
tri 17664 40268 17672 40276 ne
rect 17672 40271 17937 40276
tri 17937 40271 17945 40279 sw
rect 17672 40268 17945 40271
tri 17672 40260 17680 40268 ne
rect 17680 40263 17945 40268
tri 17945 40263 17953 40271 sw
rect 70802 40268 71000 40326
rect 17680 40260 17953 40263
tri 17680 40252 17688 40260 ne
rect 17688 40255 17953 40260
tri 17953 40255 17961 40263 sw
rect 17688 40252 17961 40255
tri 17688 40244 17696 40252 ne
rect 17696 40247 17961 40252
tri 17961 40247 17969 40255 sw
rect 17696 40244 17969 40247
tri 17696 40236 17704 40244 ne
rect 17704 40239 17969 40244
tri 17969 40239 17977 40247 sw
rect 17704 40236 17977 40239
tri 17704 40228 17712 40236 ne
rect 17712 40231 17977 40236
tri 17977 40231 17985 40239 sw
rect 17712 40228 17985 40231
tri 17712 40220 17720 40228 ne
rect 17720 40223 17985 40228
tri 17985 40223 17993 40231 sw
rect 17720 40220 17993 40223
tri 17720 40212 17728 40220 ne
rect 17728 40215 17993 40220
tri 17993 40215 18001 40223 sw
rect 70802 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17728 40212 18001 40215
tri 17728 40207 17733 40212 ne
rect 17733 40207 18001 40212
tri 18001 40207 18009 40215 sw
tri 17733 40199 17741 40207 ne
rect 17741 40204 18009 40207
rect 17741 40199 17874 40204
tri 17741 40191 17749 40199 ne
rect 17749 40191 17874 40199
tri 17749 40183 17757 40191 ne
rect 17757 40183 17874 40191
tri 17757 40175 17765 40183 ne
rect 17765 40175 17874 40183
tri 17765 40167 17773 40175 ne
rect 17773 40167 17874 40175
tri 17773 40159 17781 40167 ne
rect 17781 40159 17874 40167
tri 17781 40151 17789 40159 ne
rect 17789 40158 17874 40159
rect 17920 40199 18009 40204
tri 18009 40199 18017 40207 sw
rect 17920 40191 18017 40199
tri 18017 40191 18025 40199 sw
rect 17920 40183 18025 40191
tri 18025 40183 18033 40191 sw
rect 17920 40175 18033 40183
tri 18033 40175 18041 40183 sw
rect 17920 40167 18041 40175
tri 18041 40167 18049 40175 sw
rect 17920 40159 18049 40167
tri 18049 40159 18057 40167 sw
rect 70802 40164 71000 40222
rect 17920 40158 18057 40159
rect 17789 40151 18057 40158
tri 18057 40151 18065 40159 sw
tri 17789 40143 17797 40151 ne
rect 17797 40143 18065 40151
tri 18065 40143 18073 40151 sw
tri 17797 40140 17800 40143 ne
rect 17800 40140 18073 40143
tri 17800 40132 17808 40140 ne
rect 17808 40136 18073 40140
tri 18073 40136 18080 40143 sw
rect 17808 40132 18080 40136
tri 17808 40124 17816 40132 ne
rect 17816 40128 18080 40132
tri 18080 40128 18088 40136 sw
rect 17816 40124 18088 40128
tri 17816 40116 17824 40124 ne
rect 17824 40120 18088 40124
tri 18088 40120 18096 40128 sw
rect 17824 40116 18096 40120
tri 17824 40108 17832 40116 ne
rect 17832 40112 18096 40116
tri 18096 40112 18104 40120 sw
rect 70802 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
rect 17832 40108 18104 40112
tri 17832 40100 17840 40108 ne
rect 17840 40104 18104 40108
tri 18104 40104 18112 40112 sw
rect 17840 40100 18112 40104
tri 17840 40092 17848 40100 ne
rect 17848 40096 18112 40100
tri 18112 40096 18120 40104 sw
rect 17848 40092 18120 40096
tri 17848 40084 17856 40092 ne
rect 17856 40088 18120 40092
tri 18120 40088 18128 40096 sw
rect 17856 40084 18128 40088
tri 17856 40076 17864 40084 ne
rect 17864 40080 18128 40084
tri 18128 40080 18136 40088 sw
rect 17864 40076 18136 40080
tri 17864 40068 17872 40076 ne
rect 17872 40072 18136 40076
tri 18136 40072 18144 40080 sw
rect 17872 40068 18006 40072
tri 17872 40060 17880 40068 ne
rect 17880 40060 18006 40068
tri 17880 40052 17888 40060 ne
rect 17888 40052 18006 40060
tri 17888 40044 17896 40052 ne
rect 17896 40044 18006 40052
tri 17896 40036 17904 40044 ne
rect 17904 40036 18006 40044
tri 17904 40028 17912 40036 ne
rect 17912 40028 18006 40036
tri 17912 40025 17915 40028 ne
rect 17915 40026 18006 40028
rect 18052 40064 18144 40072
tri 18144 40064 18152 40072 sw
rect 18052 40056 18152 40064
tri 18152 40056 18160 40064 sw
rect 70802 40060 71000 40118
rect 18052 40048 18160 40056
tri 18160 40048 18168 40056 sw
rect 18052 40040 18168 40048
tri 18168 40040 18176 40048 sw
rect 18052 40032 18176 40040
tri 18176 40032 18184 40040 sw
rect 18052 40031 18184 40032
tri 18184 40031 18185 40032 sw
rect 18052 40026 18185 40031
rect 17915 40025 18185 40026
tri 17915 40017 17923 40025 ne
rect 17923 40023 18185 40025
tri 18185 40023 18193 40031 sw
rect 17923 40017 18193 40023
tri 17923 40009 17931 40017 ne
rect 17931 40015 18193 40017
tri 18193 40015 18201 40023 sw
rect 17931 40009 18201 40015
tri 17931 40001 17939 40009 ne
rect 17939 40007 18201 40009
tri 18201 40007 18209 40015 sw
rect 70802 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 17939 40001 18209 40007
tri 17939 39993 17947 40001 ne
rect 17947 39999 18209 40001
tri 18209 39999 18217 40007 sw
rect 17947 39993 18217 39999
tri 17947 39985 17955 39993 ne
rect 17955 39991 18217 39993
tri 18217 39991 18225 39999 sw
rect 17955 39985 18225 39991
tri 17955 39977 17963 39985 ne
rect 17963 39983 18225 39985
tri 18225 39983 18233 39991 sw
rect 17963 39977 18233 39983
tri 17963 39969 17971 39977 ne
rect 17971 39975 18233 39977
tri 18233 39975 18241 39983 sw
rect 17971 39969 18241 39975
tri 17971 39961 17979 39969 ne
rect 17979 39967 18241 39969
tri 18241 39967 18249 39975 sw
rect 17979 39961 18249 39967
tri 17979 39953 17987 39961 ne
rect 17987 39959 18249 39961
tri 18249 39959 18257 39967 sw
rect 17987 39953 18257 39959
tri 17987 39945 17995 39953 ne
rect 17995 39951 18257 39953
tri 18257 39951 18265 39959 sw
rect 70802 39956 71000 40014
rect 17995 39945 18265 39951
tri 17995 39937 18003 39945 ne
rect 18003 39943 18265 39945
tri 18265 39943 18273 39951 sw
rect 18003 39940 18273 39943
rect 18003 39937 18138 39940
tri 18003 39929 18011 39937 ne
rect 18011 39929 18138 39937
tri 18011 39923 18017 39929 ne
rect 18017 39923 18138 39929
tri 18017 39915 18025 39923 ne
rect 18025 39915 18138 39923
tri 18025 39907 18033 39915 ne
rect 18033 39907 18138 39915
tri 18033 39899 18041 39907 ne
rect 18041 39899 18138 39907
tri 18041 39891 18049 39899 ne
rect 18049 39894 18138 39899
rect 18184 39935 18273 39940
tri 18273 39935 18281 39943 sw
rect 18184 39927 18281 39935
tri 18281 39927 18289 39935 sw
rect 18184 39923 18289 39927
tri 18289 39923 18293 39927 sw
rect 18184 39915 18293 39923
tri 18293 39915 18301 39923 sw
rect 18184 39907 18301 39915
tri 18301 39907 18309 39915 sw
rect 70802 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 18184 39899 18309 39907
tri 18309 39899 18317 39907 sw
rect 18184 39894 18317 39899
rect 18049 39891 18317 39894
tri 18317 39891 18325 39899 sw
tri 18049 39883 18057 39891 ne
rect 18057 39883 18325 39891
tri 18325 39883 18333 39891 sw
tri 18057 39875 18065 39883 ne
rect 18065 39875 18333 39883
tri 18333 39875 18341 39883 sw
tri 18065 39867 18073 39875 ne
rect 18073 39867 18341 39875
tri 18341 39867 18349 39875 sw
tri 18073 39859 18081 39867 ne
rect 18081 39859 18349 39867
tri 18349 39859 18357 39867 sw
tri 18081 39856 18084 39859 ne
rect 18084 39856 18357 39859
tri 18084 39848 18092 39856 ne
rect 18092 39852 18357 39856
tri 18357 39852 18364 39859 sw
rect 70802 39852 71000 39910
rect 18092 39848 18364 39852
tri 18092 39840 18100 39848 ne
rect 18100 39844 18364 39848
tri 18364 39844 18372 39852 sw
rect 18100 39840 18372 39844
tri 18100 39832 18108 39840 ne
rect 18108 39836 18372 39840
tri 18372 39836 18380 39844 sw
rect 18108 39832 18380 39836
tri 18108 39824 18116 39832 ne
rect 18116 39828 18380 39832
tri 18380 39828 18388 39836 sw
rect 18116 39824 18388 39828
tri 18116 39816 18124 39824 ne
rect 18124 39820 18388 39824
tri 18388 39820 18396 39828 sw
rect 18124 39816 18396 39820
tri 18124 39808 18132 39816 ne
rect 18132 39812 18396 39816
tri 18396 39812 18404 39820 sw
rect 18132 39808 18404 39812
tri 18132 39800 18140 39808 ne
rect 18140 39800 18270 39808
tri 18140 39792 18148 39800 ne
rect 18148 39792 18270 39800
tri 18148 39784 18156 39792 ne
rect 18156 39784 18270 39792
tri 18156 39776 18164 39784 ne
rect 18164 39776 18270 39784
tri 18164 39768 18172 39776 ne
rect 18172 39768 18270 39776
tri 18172 39760 18180 39768 ne
rect 18180 39762 18270 39768
rect 18316 39804 18404 39808
tri 18404 39804 18412 39812 sw
rect 70802 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39796 18412 39804
tri 18412 39796 18420 39804 sw
rect 18316 39788 18420 39796
tri 18420 39788 18428 39796 sw
rect 18316 39780 18428 39788
tri 18428 39780 18436 39788 sw
rect 18316 39772 18436 39780
tri 18436 39772 18444 39780 sw
rect 18316 39764 18444 39772
tri 18444 39764 18452 39772 sw
rect 18316 39762 18452 39764
rect 18180 39760 18452 39762
tri 18180 39752 18188 39760 ne
rect 18188 39756 18452 39760
tri 18452 39756 18460 39764 sw
rect 18188 39755 18460 39756
tri 18460 39755 18461 39756 sw
rect 18188 39752 18461 39755
tri 18188 39751 18189 39752 ne
rect 18189 39751 18461 39752
tri 18189 39743 18197 39751 ne
rect 18197 39747 18461 39751
tri 18461 39747 18469 39755 sw
rect 70802 39748 71000 39806
rect 18197 39743 18469 39747
tri 18197 39735 18205 39743 ne
rect 18205 39739 18469 39743
tri 18469 39739 18477 39747 sw
rect 18205 39735 18477 39739
tri 18205 39727 18213 39735 ne
rect 18213 39731 18477 39735
tri 18477 39731 18485 39739 sw
rect 18213 39727 18485 39731
tri 18213 39719 18221 39727 ne
rect 18221 39723 18485 39727
tri 18485 39723 18493 39731 sw
rect 18221 39719 18493 39723
tri 18221 39711 18229 39719 ne
rect 18229 39715 18493 39719
tri 18493 39715 18501 39723 sw
rect 18229 39711 18501 39715
tri 18229 39703 18237 39711 ne
rect 18237 39707 18501 39711
tri 18501 39707 18509 39715 sw
rect 18237 39703 18509 39707
tri 18237 39695 18245 39703 ne
rect 18245 39699 18509 39703
tri 18509 39699 18517 39707 sw
rect 70802 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 18245 39695 18517 39699
tri 18245 39687 18253 39695 ne
rect 18253 39691 18517 39695
tri 18517 39691 18525 39699 sw
rect 18253 39687 18525 39691
tri 18253 39679 18261 39687 ne
rect 18261 39683 18525 39687
tri 18525 39683 18533 39691 sw
rect 18261 39679 18533 39683
tri 18261 39671 18269 39679 ne
rect 18269 39676 18533 39679
rect 18269 39671 18402 39676
tri 18269 39663 18277 39671 ne
rect 18277 39663 18402 39671
tri 18277 39655 18285 39663 ne
rect 18285 39655 18402 39663
tri 18285 39647 18293 39655 ne
rect 18293 39647 18402 39655
tri 18293 39643 18297 39647 ne
rect 18297 39643 18402 39647
tri 18297 39635 18305 39643 ne
rect 18305 39635 18402 39643
tri 18305 39627 18313 39635 ne
rect 18313 39630 18402 39635
rect 18448 39675 18533 39676
tri 18533 39675 18541 39683 sw
rect 18448 39671 18541 39675
tri 18541 39671 18545 39675 sw
rect 18448 39663 18545 39671
tri 18545 39663 18553 39671 sw
rect 18448 39655 18553 39663
tri 18553 39655 18561 39663 sw
rect 18448 39647 18561 39655
tri 18561 39647 18569 39655 sw
rect 18448 39639 18569 39647
tri 18569 39639 18577 39647 sw
rect 70802 39644 71000 39702
rect 18448 39635 18577 39639
tri 18577 39635 18581 39639 sw
rect 18448 39630 18581 39635
rect 18313 39627 18581 39630
tri 18581 39627 18589 39635 sw
tri 18313 39619 18321 39627 ne
rect 18321 39619 18589 39627
tri 18589 39619 18597 39627 sw
tri 18321 39611 18329 39619 ne
rect 18329 39611 18597 39619
tri 18597 39611 18605 39619 sw
tri 18329 39603 18337 39611 ne
rect 18337 39603 18605 39611
tri 18605 39603 18613 39611 sw
tri 18337 39595 18345 39603 ne
rect 18345 39595 18613 39603
tri 18613 39595 18621 39603 sw
rect 70802 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18345 39587 18353 39595 ne
rect 18353 39587 18621 39595
tri 18621 39587 18629 39595 sw
tri 18353 39579 18361 39587 ne
rect 18361 39579 18629 39587
tri 18629 39579 18637 39587 sw
tri 18361 39571 18369 39579 ne
rect 18369 39571 18637 39579
tri 18637 39571 18645 39579 sw
tri 18369 39563 18377 39571 ne
rect 18377 39563 18645 39571
tri 18645 39563 18653 39571 sw
tri 18377 39555 18385 39563 ne
rect 18385 39555 18653 39563
tri 18653 39555 18661 39563 sw
tri 18385 39547 18393 39555 ne
rect 18393 39547 18661 39555
tri 18661 39547 18669 39555 sw
tri 18393 39539 18401 39547 ne
rect 18401 39544 18669 39547
rect 18401 39539 18534 39544
tri 18401 39531 18409 39539 ne
rect 18409 39531 18534 39539
tri 18409 39523 18417 39531 ne
rect 18417 39523 18534 39531
tri 18417 39515 18425 39523 ne
rect 18425 39515 18534 39523
tri 18425 39513 18427 39515 ne
rect 18427 39513 18534 39515
tri 18427 39505 18435 39513 ne
rect 18435 39505 18534 39513
tri 18435 39497 18443 39505 ne
rect 18443 39498 18534 39505
rect 18580 39539 18669 39544
tri 18669 39539 18677 39547 sw
rect 70802 39540 71000 39598
rect 18580 39531 18677 39539
tri 18677 39531 18685 39539 sw
rect 18580 39523 18685 39531
tri 18685 39523 18693 39531 sw
rect 18580 39515 18693 39523
tri 18693 39515 18701 39523 sw
rect 18580 39513 18701 39515
tri 18701 39513 18703 39515 sw
rect 18580 39505 18703 39513
tri 18703 39505 18711 39513 sw
rect 18580 39498 18711 39505
rect 18443 39497 18711 39498
tri 18711 39497 18719 39505 sw
tri 18443 39489 18451 39497 ne
rect 18451 39489 18719 39497
tri 18719 39489 18727 39497 sw
rect 70802 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18451 39481 18459 39489 ne
rect 18459 39481 18727 39489
tri 18727 39481 18735 39489 sw
tri 18459 39473 18467 39481 ne
rect 18467 39473 18735 39481
tri 18735 39473 18743 39481 sw
tri 18467 39465 18475 39473 ne
rect 18475 39465 18743 39473
tri 18743 39465 18751 39473 sw
tri 18475 39457 18483 39465 ne
rect 18483 39457 18751 39465
tri 18751 39457 18759 39465 sw
tri 18483 39449 18491 39457 ne
rect 18491 39449 18759 39457
tri 18759 39449 18767 39457 sw
tri 18491 39441 18499 39449 ne
rect 18499 39441 18767 39449
tri 18767 39441 18775 39449 sw
tri 18499 39433 18507 39441 ne
rect 18507 39433 18775 39441
tri 18775 39433 18783 39441 sw
rect 70802 39436 71000 39494
tri 18507 39425 18515 39433 ne
rect 18515 39425 18783 39433
tri 18783 39425 18791 39433 sw
tri 18515 39417 18523 39425 ne
rect 18523 39417 18791 39425
tri 18791 39417 18799 39425 sw
tri 18523 39409 18531 39417 ne
rect 18531 39412 18799 39417
rect 18531 39409 18666 39412
tri 18531 39401 18539 39409 ne
rect 18539 39401 18666 39409
tri 18539 39395 18545 39401 ne
rect 18545 39395 18666 39401
tri 18545 39387 18553 39395 ne
rect 18553 39387 18666 39395
tri 18553 39379 18561 39387 ne
rect 18561 39379 18666 39387
tri 18561 39371 18569 39379 ne
rect 18569 39371 18666 39379
tri 18569 39363 18577 39371 ne
rect 18577 39366 18666 39371
rect 18712 39409 18799 39412
tri 18799 39409 18807 39417 sw
rect 18712 39401 18807 39409
tri 18807 39401 18815 39409 sw
rect 18712 39395 18815 39401
tri 18815 39395 18821 39401 sw
rect 18712 39387 18821 39395
tri 18821 39387 18829 39395 sw
rect 70802 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 18712 39379 18829 39387
tri 18829 39379 18837 39387 sw
rect 18712 39371 18837 39379
tri 18837 39371 18845 39379 sw
rect 18712 39366 18845 39371
rect 18577 39363 18845 39366
tri 18845 39363 18853 39371 sw
tri 18577 39355 18585 39363 ne
rect 18585 39355 18853 39363
tri 18853 39355 18861 39363 sw
tri 18585 39347 18593 39355 ne
rect 18593 39347 18861 39355
tri 18861 39347 18869 39355 sw
tri 18593 39339 18601 39347 ne
rect 18601 39339 18869 39347
tri 18869 39339 18877 39347 sw
tri 18601 39331 18609 39339 ne
rect 18609 39331 18877 39339
tri 18877 39331 18885 39339 sw
rect 70802 39332 71000 39390
tri 18609 39323 18617 39331 ne
rect 18617 39323 18885 39331
tri 18885 39323 18893 39331 sw
tri 18617 39315 18625 39323 ne
rect 18625 39315 18893 39323
tri 18893 39315 18901 39323 sw
tri 18625 39307 18633 39315 ne
rect 18633 39307 18901 39315
tri 18901 39307 18909 39315 sw
tri 18633 39299 18641 39307 ne
rect 18641 39299 18909 39307
tri 18909 39299 18917 39307 sw
tri 18641 39291 18649 39299 ne
rect 18649 39291 18917 39299
tri 18917 39291 18925 39299 sw
tri 18649 39283 18657 39291 ne
rect 18657 39283 18925 39291
tri 18925 39283 18933 39291 sw
rect 70802 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
tri 18657 39275 18665 39283 ne
rect 18665 39280 18933 39283
rect 18665 39275 18798 39280
tri 18665 39267 18673 39275 ne
rect 18673 39267 18798 39275
tri 18673 39259 18681 39267 ne
rect 18681 39259 18798 39267
tri 18681 39251 18689 39259 ne
rect 18689 39251 18798 39259
tri 18689 39243 18697 39251 ne
rect 18697 39243 18798 39251
tri 18697 39235 18705 39243 ne
rect 18705 39235 18798 39243
tri 18705 39227 18713 39235 ne
rect 18713 39234 18798 39235
rect 18844 39275 18933 39280
tri 18933 39275 18941 39283 sw
rect 18844 39274 18941 39275
tri 18941 39274 18942 39275 sw
rect 18844 39266 18942 39274
tri 18942 39266 18950 39274 sw
rect 18844 39258 18950 39266
tri 18950 39258 18958 39266 sw
rect 18844 39250 18958 39258
tri 18958 39250 18966 39258 sw
rect 18844 39242 18966 39250
tri 18966 39242 18974 39250 sw
rect 18844 39234 18974 39242
tri 18974 39234 18982 39242 sw
rect 18713 39227 18982 39234
tri 18713 39219 18721 39227 ne
rect 18721 39226 18982 39227
tri 18982 39226 18990 39234 sw
rect 70802 39228 71000 39286
rect 18721 39219 18990 39226
tri 18721 39211 18729 39219 ne
rect 18729 39218 18990 39219
tri 18990 39218 18998 39226 sw
rect 18729 39211 18998 39218
tri 18729 39203 18737 39211 ne
rect 18737 39210 18998 39211
tri 18998 39210 19006 39218 sw
rect 18737 39203 19006 39210
tri 18737 39195 18745 39203 ne
rect 18745 39202 19006 39203
tri 19006 39202 19014 39210 sw
rect 18745 39195 19014 39202
tri 18745 39187 18753 39195 ne
rect 18753 39194 19014 39195
tri 19014 39194 19022 39202 sw
rect 18753 39187 19022 39194
tri 18753 39179 18761 39187 ne
rect 18761 39186 19022 39187
tri 19022 39186 19030 39194 sw
rect 18761 39179 19030 39186
tri 18761 39171 18769 39179 ne
rect 18769 39178 19030 39179
tri 19030 39178 19038 39186 sw
rect 70802 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 18769 39171 19038 39178
tri 18769 39163 18777 39171 ne
rect 18777 39170 19038 39171
tri 19038 39170 19046 39178 sw
rect 18777 39167 19046 39170
tri 19046 39167 19049 39170 sw
rect 18777 39163 19049 39167
tri 18777 39159 18781 39163 ne
rect 18781 39159 19049 39163
tri 19049 39159 19057 39167 sw
tri 18781 39151 18789 39159 ne
rect 18789 39151 19057 39159
tri 19057 39151 19065 39159 sw
tri 18789 39143 18797 39151 ne
rect 18797 39148 19065 39151
rect 18797 39143 18930 39148
tri 18797 39135 18805 39143 ne
rect 18805 39135 18930 39143
tri 18805 39127 18813 39135 ne
rect 18813 39127 18930 39135
tri 18813 39119 18821 39127 ne
rect 18821 39119 18930 39127
tri 18821 39111 18829 39119 ne
rect 18829 39111 18930 39119
tri 18829 39103 18837 39111 ne
rect 18837 39103 18930 39111
tri 18837 39095 18845 39103 ne
rect 18845 39102 18930 39103
rect 18976 39143 19065 39148
tri 19065 39143 19073 39151 sw
rect 18976 39135 19073 39143
tri 19073 39135 19081 39143 sw
rect 18976 39127 19081 39135
tri 19081 39127 19089 39135 sw
rect 18976 39119 19089 39127
tri 19089 39119 19097 39127 sw
rect 70802 39124 71000 39182
rect 18976 39111 19097 39119
tri 19097 39111 19105 39119 sw
rect 18976 39103 19105 39111
tri 19105 39103 19113 39111 sw
rect 18976 39102 19113 39103
rect 18845 39095 19113 39102
tri 19113 39095 19121 39103 sw
tri 18845 39089 18851 39095 ne
rect 18851 39089 19121 39095
tri 19121 39089 19127 39095 sw
tri 18851 39081 18859 39089 ne
rect 18859 39081 19127 39089
tri 19127 39081 19135 39089 sw
tri 18859 39073 18867 39081 ne
rect 18867 39073 19135 39081
tri 19135 39073 19143 39081 sw
rect 70802 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18867 39065 18875 39073 ne
rect 18875 39065 19143 39073
tri 19143 39065 19151 39073 sw
tri 18875 39057 18883 39065 ne
rect 18883 39057 19151 39065
tri 19151 39057 19159 39065 sw
tri 18883 39049 18891 39057 ne
rect 18891 39049 19159 39057
tri 19159 39049 19167 39057 sw
tri 18891 39041 18899 39049 ne
rect 18899 39041 19167 39049
tri 19167 39041 19175 39049 sw
tri 18899 39033 18907 39041 ne
rect 18907 39033 19175 39041
tri 19175 39033 19183 39041 sw
tri 18907 39025 18915 39033 ne
rect 18915 39025 19183 39033
tri 19183 39025 19191 39033 sw
tri 18915 39017 18923 39025 ne
rect 18923 39017 19191 39025
tri 19191 39017 19199 39025 sw
rect 70802 39020 71000 39078
tri 18923 39009 18931 39017 ne
rect 18931 39016 19199 39017
rect 18931 39009 19062 39016
tri 18931 39001 18939 39009 ne
rect 18939 39001 19062 39009
tri 18939 38993 18947 39001 ne
rect 18947 38993 19062 39001
tri 18947 38985 18955 38993 ne
rect 18955 38985 19062 38993
tri 18955 38977 18963 38985 ne
rect 18963 38977 19062 38985
tri 18963 38969 18971 38977 ne
rect 18971 38970 19062 38977
rect 19108 39009 19199 39016
tri 19199 39009 19207 39017 sw
rect 19108 39001 19207 39009
tri 19207 39001 19215 39009 sw
rect 19108 38993 19215 39001
tri 19215 38993 19223 39001 sw
rect 19108 38985 19223 38993
tri 19223 38985 19231 38993 sw
rect 19108 38977 19231 38985
tri 19231 38977 19239 38985 sw
rect 19108 38970 19239 38977
rect 18971 38969 19239 38970
tri 19239 38969 19247 38977 sw
rect 70802 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
tri 18971 38961 18979 38969 ne
rect 18979 38961 19247 38969
tri 19247 38961 19255 38969 sw
tri 18979 38953 18987 38961 ne
rect 18987 38953 19255 38961
tri 19255 38953 19263 38961 sw
tri 18987 38947 18993 38953 ne
rect 18993 38947 19263 38953
tri 19263 38947 19269 38953 sw
tri 18993 38939 19001 38947 ne
rect 19001 38939 19269 38947
tri 19269 38939 19277 38947 sw
tri 19001 38931 19009 38939 ne
rect 19009 38931 19277 38939
tri 19277 38931 19285 38939 sw
tri 19009 38923 19017 38931 ne
rect 19017 38923 19285 38931
tri 19285 38923 19293 38931 sw
tri 19017 38915 19025 38923 ne
rect 19025 38915 19293 38923
tri 19293 38915 19301 38923 sw
rect 70802 38916 71000 38974
tri 19025 38907 19033 38915 ne
rect 19033 38907 19301 38915
tri 19301 38907 19309 38915 sw
tri 19033 38899 19041 38907 ne
rect 19041 38899 19309 38907
tri 19309 38899 19317 38907 sw
tri 19041 38891 19049 38899 ne
rect 19049 38891 19317 38899
tri 19317 38891 19325 38899 sw
tri 19049 38883 19057 38891 ne
rect 19057 38884 19325 38891
rect 19057 38883 19194 38884
tri 19057 38875 19065 38883 ne
rect 19065 38875 19194 38883
tri 19065 38867 19073 38875 ne
rect 19073 38867 19194 38875
tri 19073 38859 19081 38867 ne
rect 19081 38859 19194 38867
tri 19081 38851 19089 38859 ne
rect 19089 38851 19194 38859
tri 19089 38843 19097 38851 ne
rect 19097 38843 19194 38851
tri 19097 38835 19105 38843 ne
rect 19105 38838 19194 38843
rect 19240 38883 19325 38884
tri 19325 38883 19333 38891 sw
rect 19240 38875 19333 38883
tri 19333 38875 19341 38883 sw
rect 19240 38867 19341 38875
tri 19341 38867 19349 38875 sw
rect 70802 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38859 19349 38867
tri 19349 38859 19357 38867 sw
rect 19240 38851 19357 38859
tri 19357 38851 19365 38859 sw
rect 19240 38843 19365 38851
tri 19365 38843 19373 38851 sw
rect 19240 38838 19373 38843
rect 19105 38835 19373 38838
tri 19373 38835 19381 38843 sw
tri 19105 38827 19113 38835 ne
rect 19113 38827 19381 38835
tri 19381 38827 19389 38835 sw
tri 19113 38819 19121 38827 ne
rect 19121 38819 19389 38827
tri 19389 38819 19397 38827 sw
tri 19121 38811 19129 38819 ne
rect 19129 38811 19397 38819
tri 19397 38811 19405 38819 sw
rect 70802 38812 71000 38870
tri 19129 38805 19135 38811 ne
rect 19135 38805 19405 38811
tri 19405 38805 19411 38811 sw
tri 19135 38797 19143 38805 ne
rect 19143 38797 19411 38805
tri 19411 38797 19419 38805 sw
tri 19143 38789 19151 38797 ne
rect 19151 38789 19419 38797
tri 19419 38789 19427 38797 sw
tri 19151 38781 19159 38789 ne
rect 19159 38781 19427 38789
tri 19427 38781 19435 38789 sw
tri 19159 38773 19167 38781 ne
rect 19167 38773 19435 38781
tri 19435 38773 19443 38781 sw
tri 19167 38765 19175 38773 ne
rect 19175 38765 19443 38773
tri 19443 38765 19451 38773 sw
rect 70802 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19175 38757 19183 38765 ne
rect 19183 38757 19451 38765
tri 19451 38757 19459 38765 sw
tri 19183 38749 19191 38757 ne
rect 19191 38752 19459 38757
rect 19191 38749 19326 38752
tri 19191 38741 19199 38749 ne
rect 19199 38741 19326 38749
tri 19199 38733 19207 38741 ne
rect 19207 38733 19326 38741
tri 19207 38725 19215 38733 ne
rect 19215 38725 19326 38733
tri 19215 38717 19223 38725 ne
rect 19223 38717 19326 38725
tri 19223 38709 19231 38717 ne
rect 19231 38709 19326 38717
tri 19231 38701 19239 38709 ne
rect 19239 38706 19326 38709
rect 19372 38749 19459 38752
tri 19459 38749 19467 38757 sw
rect 19372 38741 19467 38749
tri 19467 38741 19475 38749 sw
rect 19372 38733 19475 38741
tri 19475 38733 19483 38741 sw
rect 19372 38725 19483 38733
tri 19483 38725 19491 38733 sw
rect 19372 38717 19491 38725
tri 19491 38717 19499 38725 sw
rect 19372 38709 19499 38717
tri 19499 38709 19507 38717 sw
rect 19372 38706 19507 38709
rect 19239 38701 19507 38706
tri 19507 38701 19515 38709 sw
rect 70802 38708 71000 38766
tri 19239 38695 19245 38701 ne
rect 19245 38695 19515 38701
tri 19515 38695 19521 38701 sw
tri 19245 38687 19253 38695 ne
rect 19253 38687 19521 38695
tri 19521 38687 19529 38695 sw
tri 19253 38679 19261 38687 ne
rect 19261 38679 19529 38687
tri 19529 38679 19537 38687 sw
tri 19261 38671 19269 38679 ne
rect 19269 38671 19537 38679
tri 19537 38671 19545 38679 sw
tri 19269 38663 19277 38671 ne
rect 19277 38663 19545 38671
tri 19545 38663 19553 38671 sw
tri 19277 38655 19285 38663 ne
rect 19285 38655 19553 38663
tri 19553 38655 19561 38663 sw
rect 70802 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19285 38647 19293 38655 ne
rect 19293 38647 19561 38655
tri 19561 38647 19569 38655 sw
tri 19293 38639 19301 38647 ne
rect 19301 38639 19569 38647
tri 19569 38639 19577 38647 sw
tri 19301 38631 19309 38639 ne
rect 19309 38631 19577 38639
tri 19577 38631 19585 38639 sw
tri 19309 38623 19317 38631 ne
rect 19317 38623 19585 38631
tri 19585 38623 19593 38631 sw
tri 19317 38615 19325 38623 ne
rect 19325 38620 19593 38623
rect 19325 38615 19458 38620
tri 19325 38607 19333 38615 ne
rect 19333 38607 19458 38615
tri 19333 38599 19341 38607 ne
rect 19341 38599 19458 38607
tri 19341 38591 19349 38599 ne
rect 19349 38591 19458 38599
tri 19349 38583 19357 38591 ne
rect 19357 38583 19458 38591
tri 19357 38575 19365 38583 ne
rect 19365 38575 19458 38583
tri 19365 38567 19373 38575 ne
rect 19373 38574 19458 38575
rect 19504 38615 19593 38620
tri 19593 38615 19601 38623 sw
rect 19504 38607 19601 38615
tri 19601 38607 19609 38615 sw
rect 19504 38599 19609 38607
tri 19609 38599 19617 38607 sw
rect 70802 38604 71000 38662
rect 19504 38591 19617 38599
tri 19617 38591 19625 38599 sw
rect 19504 38583 19625 38591
tri 19625 38583 19633 38591 sw
rect 19504 38575 19633 38583
tri 19633 38575 19641 38583 sw
rect 19504 38574 19641 38575
rect 19373 38567 19641 38574
tri 19641 38567 19649 38575 sw
tri 19373 38559 19381 38567 ne
rect 19381 38559 19649 38567
tri 19649 38559 19657 38567 sw
tri 19381 38553 19387 38559 ne
rect 19387 38553 19657 38559
tri 19657 38553 19663 38559 sw
rect 70802 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
tri 19387 38545 19395 38553 ne
rect 19395 38545 19663 38553
tri 19663 38545 19671 38553 sw
tri 19395 38537 19403 38545 ne
rect 19403 38537 19671 38545
tri 19671 38537 19679 38545 sw
tri 19403 38529 19411 38537 ne
rect 19411 38529 19679 38537
tri 19679 38529 19687 38537 sw
tri 19411 38521 19419 38529 ne
rect 19419 38521 19687 38529
tri 19687 38521 19695 38529 sw
tri 19419 38513 19427 38521 ne
rect 19427 38513 19695 38521
tri 19695 38513 19703 38521 sw
tri 19427 38505 19435 38513 ne
rect 19435 38505 19703 38513
tri 19703 38505 19711 38513 sw
tri 19435 38497 19443 38505 ne
rect 19443 38497 19711 38505
tri 19711 38497 19719 38505 sw
rect 70802 38500 71000 38558
tri 19443 38489 19451 38497 ne
rect 19451 38489 19719 38497
tri 19719 38489 19727 38497 sw
tri 19451 38481 19459 38489 ne
rect 19459 38488 19727 38489
rect 19459 38481 19590 38488
tri 19459 38473 19467 38481 ne
rect 19467 38473 19590 38481
tri 19467 38465 19475 38473 ne
rect 19475 38465 19590 38473
tri 19475 38457 19483 38465 ne
rect 19483 38457 19590 38465
tri 19483 38449 19491 38457 ne
rect 19491 38449 19590 38457
tri 19491 38441 19499 38449 ne
rect 19499 38442 19590 38449
rect 19636 38481 19727 38488
tri 19727 38481 19735 38489 sw
rect 19636 38473 19735 38481
tri 19735 38473 19743 38481 sw
rect 19636 38465 19743 38473
tri 19743 38465 19751 38473 sw
rect 19636 38457 19751 38465
tri 19751 38457 19759 38465 sw
rect 19636 38449 19759 38457
tri 19759 38449 19767 38457 sw
rect 70802 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19767 38449
rect 19499 38441 19767 38442
tri 19767 38441 19775 38449 sw
tri 19499 38433 19507 38441 ne
rect 19507 38433 19775 38441
tri 19775 38433 19783 38441 sw
tri 19507 38425 19515 38433 ne
rect 19515 38425 19783 38433
tri 19783 38425 19791 38433 sw
tri 19515 38417 19523 38425 ne
rect 19523 38417 19791 38425
tri 19791 38417 19799 38425 sw
tri 19523 38411 19529 38417 ne
rect 19529 38411 19799 38417
tri 19799 38411 19805 38417 sw
tri 19529 38403 19537 38411 ne
rect 19537 38403 19805 38411
tri 19805 38403 19813 38411 sw
tri 19537 38395 19545 38403 ne
rect 19545 38395 19813 38403
tri 19813 38395 19821 38403 sw
rect 70802 38396 71000 38454
tri 19545 38387 19553 38395 ne
rect 19553 38387 19821 38395
tri 19821 38387 19829 38395 sw
tri 19553 38379 19561 38387 ne
rect 19561 38379 19829 38387
tri 19829 38379 19837 38387 sw
tri 19561 38371 19569 38379 ne
rect 19569 38371 19837 38379
tri 19837 38371 19845 38379 sw
tri 19569 38363 19577 38371 ne
rect 19577 38363 19845 38371
tri 19845 38363 19853 38371 sw
tri 19577 38355 19585 38363 ne
rect 19585 38356 19853 38363
rect 19585 38355 19722 38356
tri 19585 38347 19593 38355 ne
rect 19593 38347 19722 38355
tri 19593 38339 19601 38347 ne
rect 19601 38339 19722 38347
tri 19601 38331 19609 38339 ne
rect 19609 38331 19722 38339
tri 19609 38323 19617 38331 ne
rect 19617 38323 19722 38331
tri 19617 38315 19625 38323 ne
rect 19625 38315 19722 38323
tri 19625 38307 19633 38315 ne
rect 19633 38310 19722 38315
rect 19768 38355 19853 38356
tri 19853 38355 19861 38363 sw
rect 19768 38347 19861 38355
tri 19861 38347 19869 38355 sw
rect 70802 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 19768 38339 19869 38347
tri 19869 38339 19877 38347 sw
rect 19768 38331 19877 38339
tri 19877 38331 19885 38339 sw
rect 19768 38323 19885 38331
tri 19885 38323 19893 38331 sw
rect 19768 38315 19893 38323
tri 19893 38315 19901 38323 sw
rect 19768 38310 19901 38315
rect 19633 38307 19901 38310
tri 19901 38307 19909 38315 sw
tri 19633 38299 19641 38307 ne
rect 19641 38299 19909 38307
tri 19909 38299 19917 38307 sw
tri 19641 38291 19649 38299 ne
rect 19649 38291 19917 38299
tri 19917 38291 19925 38299 sw
rect 70802 38292 71000 38350
tri 19649 38283 19657 38291 ne
rect 19657 38290 19925 38291
tri 19925 38290 19926 38291 sw
rect 19657 38283 19926 38290
tri 19657 38275 19665 38283 ne
rect 19665 38282 19926 38283
tri 19926 38282 19934 38290 sw
rect 19665 38275 19934 38282
tri 19665 38274 19666 38275 ne
rect 19666 38274 19934 38275
tri 19934 38274 19942 38282 sw
tri 19666 38266 19674 38274 ne
rect 19674 38266 19942 38274
tri 19942 38266 19950 38274 sw
tri 19674 38258 19682 38266 ne
rect 19682 38258 19950 38266
tri 19950 38258 19958 38266 sw
tri 19682 38250 19690 38258 ne
rect 19690 38250 19958 38258
tri 19958 38250 19966 38258 sw
tri 19690 38242 19698 38250 ne
rect 19698 38242 19966 38250
tri 19966 38242 19974 38250 sw
rect 70802 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
tri 19698 38234 19706 38242 ne
rect 19706 38234 19974 38242
tri 19974 38234 19982 38242 sw
tri 19706 38226 19714 38234 ne
rect 19714 38226 19982 38234
tri 19982 38226 19990 38234 sw
tri 19714 38218 19722 38226 ne
rect 19722 38224 19990 38226
rect 19722 38218 19854 38224
tri 19722 38210 19730 38218 ne
rect 19730 38210 19854 38218
tri 19730 38202 19738 38210 ne
rect 19738 38202 19854 38210
tri 19738 38194 19746 38202 ne
rect 19746 38194 19854 38202
tri 19746 38186 19754 38194 ne
rect 19754 38186 19854 38194
tri 19754 38178 19762 38186 ne
rect 19762 38178 19854 38186
rect 19900 38218 19990 38224
tri 19990 38218 19998 38226 sw
rect 19900 38210 19998 38218
tri 19998 38210 20006 38218 sw
rect 19900 38202 20006 38210
tri 20006 38202 20014 38210 sw
rect 19900 38194 20014 38202
tri 20014 38194 20022 38202 sw
rect 19900 38186 20022 38194
tri 20022 38186 20030 38194 sw
rect 70802 38188 71000 38246
rect 19900 38183 20030 38186
tri 20030 38183 20033 38186 sw
rect 19900 38178 20033 38183
tri 19762 38170 19770 38178 ne
rect 19770 38175 20033 38178
tri 20033 38175 20041 38183 sw
rect 19770 38170 20041 38175
tri 19770 38162 19778 38170 ne
rect 19778 38167 20041 38170
tri 20041 38167 20049 38175 sw
rect 19778 38162 20049 38167
tri 19778 38159 19781 38162 ne
rect 19781 38159 20049 38162
tri 20049 38159 20057 38167 sw
tri 19781 38151 19789 38159 ne
rect 19789 38151 20057 38159
tri 20057 38151 20065 38159 sw
tri 19789 38143 19797 38151 ne
rect 19797 38143 20065 38151
tri 20065 38143 20073 38151 sw
tri 19797 38135 19805 38143 ne
rect 19805 38135 20073 38143
tri 20073 38135 20081 38143 sw
rect 70802 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
tri 19805 38127 19813 38135 ne
rect 19813 38127 20081 38135
tri 20081 38127 20089 38135 sw
tri 19813 38119 19821 38127 ne
rect 19821 38119 20089 38127
tri 20089 38119 20097 38127 sw
tri 19821 38111 19829 38119 ne
rect 19829 38111 20097 38119
tri 20097 38111 20105 38119 sw
tri 19829 38103 19837 38111 ne
rect 19837 38103 20105 38111
tri 20105 38103 20113 38111 sw
tri 19837 38095 19845 38103 ne
rect 19845 38095 20113 38103
tri 20113 38095 20121 38103 sw
tri 19845 38087 19853 38095 ne
rect 19853 38092 20121 38095
rect 19853 38087 19986 38092
tri 19853 38079 19861 38087 ne
rect 19861 38079 19986 38087
tri 19861 38071 19869 38079 ne
rect 19869 38071 19986 38079
tri 19869 38063 19877 38071 ne
rect 19877 38063 19986 38071
tri 19877 38055 19885 38063 ne
rect 19885 38055 19986 38063
tri 19885 38047 19893 38055 ne
rect 19893 38047 19986 38055
tri 19893 38039 19901 38047 ne
rect 19901 38046 19986 38047
rect 20032 38087 20121 38092
tri 20121 38087 20129 38095 sw
rect 20032 38079 20129 38087
tri 20129 38079 20137 38087 sw
rect 70802 38084 71000 38142
rect 20032 38071 20137 38079
tri 20137 38071 20145 38079 sw
rect 20032 38063 20145 38071
tri 20145 38063 20153 38071 sw
rect 20032 38055 20153 38063
tri 20153 38055 20161 38063 sw
rect 20032 38047 20161 38055
tri 20161 38047 20169 38055 sw
rect 20032 38046 20169 38047
tri 20169 38046 20170 38047 sw
rect 19901 38039 20170 38046
tri 19901 38038 19902 38039 ne
rect 19902 38038 20170 38039
tri 20170 38038 20178 38046 sw
rect 70802 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
tri 19902 38030 19910 38038 ne
rect 19910 38030 20178 38038
tri 20178 38030 20186 38038 sw
tri 19910 38022 19918 38030 ne
rect 19918 38022 20186 38030
tri 20186 38022 20194 38030 sw
tri 19918 38014 19926 38022 ne
rect 19926 38014 20194 38022
tri 20194 38014 20202 38022 sw
tri 19926 38006 19934 38014 ne
rect 19934 38006 20202 38014
tri 20202 38006 20210 38014 sw
tri 19934 37998 19942 38006 ne
rect 19942 37998 20210 38006
tri 20210 37998 20218 38006 sw
tri 19942 37990 19950 37998 ne
rect 19950 37990 20218 37998
tri 20218 37990 20226 37998 sw
tri 19950 37982 19958 37990 ne
rect 19958 37982 20226 37990
tri 20226 37982 20234 37990 sw
tri 19958 37974 19966 37982 ne
rect 19966 37974 20234 37982
tri 20234 37974 20242 37982 sw
rect 70802 37980 71000 38038
tri 19966 37966 19974 37974 ne
rect 19974 37966 20242 37974
tri 20242 37966 20250 37974 sw
tri 19974 37958 19982 37966 ne
rect 19982 37960 20250 37966
rect 19982 37958 20118 37960
tri 19982 37950 19990 37958 ne
rect 19990 37950 20118 37958
tri 19990 37942 19998 37950 ne
rect 19998 37942 20118 37950
tri 19998 37934 20006 37942 ne
rect 20006 37934 20118 37942
tri 20006 37926 20014 37934 ne
rect 20014 37926 20118 37934
tri 20014 37918 20022 37926 ne
rect 20022 37918 20118 37926
tri 20022 37911 20029 37918 ne
rect 20029 37914 20118 37918
rect 20164 37958 20250 37960
tri 20250 37958 20258 37966 sw
rect 20164 37950 20258 37958
tri 20258 37950 20266 37958 sw
rect 20164 37942 20266 37950
tri 20266 37942 20274 37950 sw
rect 20164 37934 20274 37942
tri 20274 37934 20282 37942 sw
rect 70802 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 20164 37927 20282 37934
tri 20282 37927 20289 37934 sw
rect 20164 37919 20289 37927
tri 20289 37919 20297 37927 sw
rect 20164 37914 20297 37919
rect 20029 37911 20297 37914
tri 20297 37911 20305 37919 sw
tri 20029 37903 20037 37911 ne
rect 20037 37903 20305 37911
tri 20305 37903 20313 37911 sw
tri 20037 37895 20045 37903 ne
rect 20045 37895 20313 37903
tri 20313 37895 20321 37903 sw
tri 20045 37887 20053 37895 ne
rect 20053 37887 20321 37895
tri 20321 37887 20329 37895 sw
tri 20053 37879 20061 37887 ne
rect 20061 37879 20329 37887
tri 20329 37879 20337 37887 sw
tri 20061 37871 20069 37879 ne
rect 20069 37871 20337 37879
tri 20337 37871 20345 37879 sw
rect 70802 37876 71000 37934
tri 20069 37863 20077 37871 ne
rect 20077 37863 20345 37871
tri 20345 37863 20353 37871 sw
tri 20077 37855 20085 37863 ne
rect 20085 37855 20353 37863
tri 20353 37855 20361 37863 sw
tri 20085 37847 20093 37855 ne
rect 20093 37847 20361 37855
tri 20361 37847 20369 37855 sw
tri 20093 37839 20101 37847 ne
rect 20101 37839 20369 37847
tri 20369 37839 20377 37847 sw
tri 20101 37835 20105 37839 ne
rect 20105 37835 20377 37839
tri 20377 37835 20381 37839 sw
tri 20105 37827 20113 37835 ne
rect 20113 37828 20381 37835
rect 20113 37827 20250 37828
tri 20113 37819 20121 37827 ne
rect 20121 37819 20250 37827
tri 20121 37811 20129 37819 ne
rect 20129 37811 20250 37819
tri 20129 37803 20137 37811 ne
rect 20137 37803 20250 37811
tri 20137 37795 20145 37803 ne
rect 20145 37795 20250 37803
tri 20145 37787 20153 37795 ne
rect 20153 37787 20250 37795
tri 20153 37779 20161 37787 ne
rect 20161 37782 20250 37787
rect 20296 37827 20381 37828
tri 20381 37827 20389 37835 sw
rect 70802 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 20296 37819 20389 37827
tri 20389 37819 20397 37827 sw
rect 20296 37811 20397 37819
tri 20397 37811 20405 37819 sw
rect 20296 37803 20405 37811
tri 20405 37803 20413 37811 sw
rect 20296 37795 20413 37803
tri 20413 37795 20421 37803 sw
rect 20296 37787 20421 37795
tri 20421 37787 20429 37795 sw
rect 20296 37782 20429 37787
rect 20161 37779 20429 37782
tri 20429 37779 20437 37787 sw
tri 20161 37771 20169 37779 ne
rect 20169 37771 20437 37779
tri 20437 37771 20445 37779 sw
rect 70802 37772 71000 37830
tri 20169 37763 20177 37771 ne
rect 20177 37763 20445 37771
tri 20445 37763 20453 37771 sw
tri 20177 37755 20185 37763 ne
rect 20185 37755 20453 37763
tri 20453 37755 20461 37763 sw
tri 20185 37747 20193 37755 ne
rect 20193 37747 20461 37755
tri 20461 37747 20469 37755 sw
tri 20193 37739 20201 37747 ne
rect 20201 37739 20469 37747
tri 20469 37739 20477 37747 sw
tri 20201 37731 20209 37739 ne
rect 20209 37731 20477 37739
tri 20477 37731 20485 37739 sw
tri 20209 37723 20217 37731 ne
rect 20217 37723 20485 37731
tri 20485 37723 20493 37731 sw
rect 70802 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
tri 20217 37715 20225 37723 ne
rect 20225 37715 20493 37723
tri 20493 37715 20501 37723 sw
tri 20225 37707 20233 37715 ne
rect 20233 37707 20501 37715
tri 20501 37707 20509 37715 sw
tri 20233 37699 20241 37707 ne
rect 20241 37699 20509 37707
tri 20509 37699 20517 37707 sw
tri 20241 37695 20245 37699 ne
rect 20245 37696 20517 37699
rect 20245 37695 20382 37696
tri 20245 37687 20253 37695 ne
rect 20253 37687 20382 37695
tri 20253 37679 20261 37687 ne
rect 20261 37679 20382 37687
tri 20261 37671 20269 37679 ne
rect 20269 37671 20382 37679
tri 20269 37663 20277 37671 ne
rect 20277 37663 20382 37671
tri 20277 37655 20285 37663 ne
rect 20285 37655 20382 37663
tri 20285 37647 20293 37655 ne
rect 20293 37650 20382 37655
rect 20428 37691 20517 37696
tri 20517 37691 20525 37699 sw
rect 20428 37683 20525 37691
tri 20525 37683 20533 37691 sw
rect 20428 37675 20533 37683
tri 20533 37675 20541 37683 sw
rect 20428 37667 20541 37675
tri 20541 37667 20549 37675 sw
rect 70802 37668 71000 37726
rect 20428 37659 20549 37667
tri 20549 37659 20557 37667 sw
rect 20428 37651 20557 37659
tri 20557 37651 20565 37659 sw
rect 20428 37650 20565 37651
rect 20293 37647 20565 37650
tri 20293 37639 20301 37647 ne
rect 20301 37643 20565 37647
tri 20565 37643 20573 37651 sw
rect 20301 37639 20573 37643
tri 20301 37631 20309 37639 ne
rect 20309 37635 20573 37639
tri 20573 37635 20581 37643 sw
rect 20309 37631 20581 37635
tri 20309 37623 20317 37631 ne
rect 20317 37627 20581 37631
tri 20581 37627 20589 37635 sw
rect 20317 37623 20589 37627
tri 20317 37615 20325 37623 ne
rect 20325 37619 20589 37623
tri 20589 37619 20597 37627 sw
rect 70802 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
rect 20325 37615 20597 37619
tri 20325 37607 20333 37615 ne
rect 20333 37611 20597 37615
tri 20597 37611 20605 37619 sw
rect 20333 37607 20605 37611
tri 20333 37599 20341 37607 ne
rect 20341 37603 20605 37607
tri 20605 37603 20613 37611 sw
rect 20341 37599 20613 37603
tri 20341 37591 20349 37599 ne
rect 20349 37595 20613 37599
tri 20613 37595 20621 37603 sw
rect 20349 37591 20621 37595
tri 20349 37587 20353 37591 ne
rect 20353 37587 20621 37591
tri 20621 37587 20629 37595 sw
tri 20353 37583 20357 37587 ne
rect 20357 37583 20629 37587
tri 20629 37583 20633 37587 sw
tri 20357 37575 20365 37583 ne
rect 20365 37575 20633 37583
tri 20633 37575 20641 37583 sw
tri 20365 37567 20373 37575 ne
rect 20373 37567 20641 37575
tri 20641 37567 20649 37575 sw
tri 20373 37559 20381 37567 ne
rect 20381 37564 20649 37567
rect 20381 37559 20514 37564
tri 20381 37551 20389 37559 ne
rect 20389 37551 20514 37559
tri 20389 37543 20397 37551 ne
rect 20397 37543 20514 37551
tri 20397 37535 20405 37543 ne
rect 20405 37535 20514 37543
tri 20405 37527 20413 37535 ne
rect 20413 37527 20514 37535
tri 20413 37519 20421 37527 ne
rect 20421 37519 20514 37527
tri 20421 37511 20429 37519 ne
rect 20429 37518 20514 37519
rect 20560 37559 20649 37564
tri 20649 37559 20657 37567 sw
rect 70802 37564 71000 37622
rect 20560 37551 20657 37559
tri 20657 37551 20665 37559 sw
rect 20560 37543 20665 37551
tri 20665 37543 20673 37551 sw
rect 20560 37535 20673 37543
tri 20673 37535 20681 37543 sw
rect 20560 37527 20681 37535
tri 20681 37527 20689 37535 sw
rect 20560 37523 20689 37527
tri 20689 37523 20693 37527 sw
rect 20560 37518 20693 37523
rect 20429 37515 20693 37518
tri 20693 37515 20701 37523 sw
rect 70802 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 20429 37511 20701 37515
tri 20429 37503 20437 37511 ne
rect 20437 37507 20701 37511
tri 20701 37507 20709 37515 sw
rect 20437 37503 20709 37507
tri 20437 37498 20442 37503 ne
rect 20442 37499 20709 37503
tri 20709 37499 20717 37507 sw
rect 20442 37498 20717 37499
tri 20442 37490 20450 37498 ne
rect 20450 37491 20717 37498
tri 20717 37491 20725 37499 sw
rect 20450 37490 20725 37491
tri 20450 37482 20458 37490 ne
rect 20458 37483 20725 37490
tri 20725 37483 20733 37491 sw
rect 20458 37482 20733 37483
tri 20458 37474 20466 37482 ne
rect 20466 37475 20733 37482
tri 20733 37475 20741 37483 sw
rect 20466 37474 20741 37475
tri 20466 37466 20474 37474 ne
rect 20474 37467 20741 37474
tri 20741 37467 20749 37475 sw
rect 20474 37466 20749 37467
tri 20474 37458 20482 37466 ne
rect 20482 37459 20749 37466
tri 20749 37459 20757 37467 sw
rect 70802 37460 71000 37518
rect 20482 37458 20757 37459
tri 20482 37450 20490 37458 ne
rect 20490 37451 20757 37458
tri 20757 37451 20765 37459 sw
rect 20490 37450 20765 37451
tri 20490 37442 20498 37450 ne
rect 20498 37443 20765 37450
tri 20765 37443 20773 37451 sw
rect 20498 37442 20773 37443
tri 20498 37434 20506 37442 ne
rect 20506 37435 20773 37442
tri 20773 37435 20781 37443 sw
rect 20506 37434 20781 37435
tri 20506 37426 20514 37434 ne
rect 20514 37432 20781 37434
rect 20514 37426 20646 37432
tri 20514 37418 20522 37426 ne
rect 20522 37418 20646 37426
tri 20522 37410 20530 37418 ne
rect 20530 37410 20646 37418
tri 20530 37402 20538 37410 ne
rect 20538 37402 20646 37410
tri 20538 37394 20546 37402 ne
rect 20546 37394 20646 37402
tri 20546 37386 20554 37394 ne
rect 20554 37386 20646 37394
rect 20692 37427 20781 37432
tri 20781 37427 20789 37435 sw
rect 20692 37419 20789 37427
tri 20789 37419 20797 37427 sw
rect 20692 37411 20797 37419
tri 20797 37411 20805 37419 sw
rect 70802 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 20692 37403 20805 37411
tri 20805 37403 20813 37411 sw
rect 20692 37395 20813 37403
tri 20813 37395 20821 37403 sw
rect 20692 37391 20821 37395
tri 20821 37391 20825 37395 sw
rect 20692 37386 20825 37391
tri 20554 37378 20562 37386 ne
rect 20562 37383 20825 37386
tri 20825 37383 20833 37391 sw
rect 20562 37378 20833 37383
tri 20562 37370 20570 37378 ne
rect 20570 37375 20833 37378
tri 20833 37375 20841 37383 sw
rect 20570 37370 20841 37375
tri 20570 37362 20578 37370 ne
rect 20578 37367 20841 37370
tri 20841 37367 20849 37375 sw
rect 20578 37362 20849 37367
tri 20578 37355 20585 37362 ne
rect 20585 37359 20849 37362
tri 20849 37359 20857 37367 sw
rect 20585 37355 20857 37359
tri 20585 37347 20593 37355 ne
rect 20593 37351 20857 37355
tri 20857 37351 20865 37359 sw
rect 70802 37356 71000 37414
rect 20593 37347 20865 37351
tri 20593 37339 20601 37347 ne
rect 20601 37343 20865 37347
tri 20865 37343 20873 37351 sw
rect 20601 37339 20873 37343
tri 20601 37331 20609 37339 ne
rect 20609 37335 20873 37339
tri 20873 37335 20881 37343 sw
rect 20609 37331 20881 37335
tri 20609 37323 20617 37331 ne
rect 20617 37327 20881 37331
tri 20881 37327 20889 37335 sw
rect 20617 37323 20889 37327
tri 20617 37315 20625 37323 ne
rect 20625 37319 20889 37323
tri 20889 37319 20897 37327 sw
rect 20625 37315 20897 37319
tri 20625 37307 20633 37315 ne
rect 20633 37311 20897 37315
tri 20897 37311 20905 37319 sw
rect 20633 37307 20905 37311
tri 20633 37299 20641 37307 ne
rect 20641 37303 20905 37307
tri 20905 37303 20913 37311 sw
rect 70802 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 20641 37300 20913 37303
rect 20641 37299 20778 37300
tri 20641 37295 20645 37299 ne
rect 20645 37295 20778 37299
tri 20645 37291 20649 37295 ne
rect 20649 37291 20778 37295
tri 20649 37283 20657 37291 ne
rect 20657 37283 20778 37291
tri 20657 37275 20665 37283 ne
rect 20665 37275 20778 37283
tri 20665 37267 20673 37275 ne
rect 20673 37267 20778 37275
tri 20673 37259 20681 37267 ne
rect 20681 37259 20778 37267
tri 20681 37251 20689 37259 ne
rect 20689 37254 20778 37259
rect 20824 37299 20913 37300
tri 20913 37299 20917 37303 sw
rect 20824 37291 20917 37299
tri 20917 37291 20925 37299 sw
rect 20824 37283 20925 37291
tri 20925 37283 20933 37291 sw
rect 20824 37275 20933 37283
tri 20933 37275 20941 37283 sw
rect 20824 37267 20941 37275
tri 20941 37267 20949 37275 sw
rect 20824 37259 20949 37267
tri 20949 37259 20957 37267 sw
rect 20824 37254 20957 37259
rect 20689 37251 20957 37254
tri 20957 37251 20965 37259 sw
rect 70802 37252 71000 37310
tri 20689 37243 20697 37251 ne
rect 20697 37243 20965 37251
tri 20965 37243 20973 37251 sw
tri 20697 37235 20705 37243 ne
rect 20705 37235 20973 37243
tri 20973 37235 20981 37243 sw
tri 20705 37227 20713 37235 ne
rect 20713 37227 20981 37235
tri 20981 37227 20989 37235 sw
tri 20713 37219 20721 37227 ne
rect 20721 37219 20989 37227
tri 20989 37219 20997 37227 sw
tri 20721 37211 20729 37219 ne
rect 20729 37211 20997 37219
tri 20997 37211 21005 37219 sw
tri 20729 37203 20737 37211 ne
rect 20737 37203 21005 37211
tri 21005 37203 21013 37211 sw
rect 70802 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
tri 20737 37195 20745 37203 ne
rect 20745 37195 21013 37203
tri 21013 37195 21021 37203 sw
tri 20745 37187 20753 37195 ne
rect 20753 37187 21021 37195
tri 21021 37187 21029 37195 sw
tri 20753 37179 20761 37187 ne
rect 20761 37179 21029 37187
tri 21029 37179 21037 37187 sw
tri 20761 37171 20769 37179 ne
rect 20769 37176 21037 37179
tri 21037 37176 21040 37179 sw
rect 20769 37171 21040 37176
tri 20769 37163 20777 37171 ne
rect 20777 37168 21040 37171
tri 21040 37168 21048 37176 sw
rect 20777 37163 20910 37168
tri 20777 37159 20781 37163 ne
rect 20781 37159 20910 37163
tri 20781 37151 20789 37159 ne
rect 20789 37151 20910 37159
tri 20789 37143 20797 37151 ne
rect 20797 37143 20910 37151
tri 20797 37135 20805 37143 ne
rect 20805 37135 20910 37143
tri 20805 37127 20813 37135 ne
rect 20813 37127 20910 37135
tri 20813 37119 20821 37127 ne
rect 20821 37122 20910 37127
rect 20956 37160 21048 37168
tri 21048 37160 21056 37168 sw
rect 20956 37152 21056 37160
tri 21056 37152 21064 37160 sw
rect 20956 37144 21064 37152
tri 21064 37144 21072 37152 sw
rect 70802 37148 71000 37206
rect 20956 37136 21072 37144
tri 21072 37136 21080 37144 sw
rect 20956 37128 21080 37136
tri 21080 37128 21088 37136 sw
rect 20956 37122 21088 37128
rect 20821 37120 21088 37122
tri 21088 37120 21096 37128 sw
rect 20821 37119 21096 37120
tri 20821 37111 20829 37119 ne
rect 20829 37112 21096 37119
tri 21096 37112 21104 37120 sw
rect 20829 37111 21104 37112
tri 20829 37103 20837 37111 ne
rect 20837 37104 21104 37111
tri 21104 37104 21112 37112 sw
rect 20837 37103 21112 37104
tri 20837 37095 20845 37103 ne
rect 20845 37096 21112 37103
tri 21112 37096 21120 37104 sw
rect 70802 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
rect 20845 37095 21120 37096
tri 20845 37087 20853 37095 ne
rect 20853 37088 21120 37095
tri 21120 37088 21128 37096 sw
rect 20853 37087 21128 37088
tri 20853 37079 20861 37087 ne
rect 20861 37080 21128 37087
tri 21128 37080 21136 37088 sw
rect 20861 37079 21136 37080
tri 20861 37071 20869 37079 ne
rect 20869 37072 21136 37079
tri 21136 37072 21144 37080 sw
rect 20869 37071 21144 37072
tri 20869 37063 20877 37071 ne
rect 20877 37064 21144 37071
tri 21144 37064 21152 37072 sw
rect 20877 37063 21152 37064
tri 21152 37063 21153 37064 sw
tri 20877 37055 20885 37063 ne
rect 20885 37055 21153 37063
tri 21153 37055 21161 37063 sw
tri 20885 37047 20893 37055 ne
rect 20893 37047 21161 37055
tri 21161 37047 21169 37055 sw
tri 20893 37039 20901 37047 ne
rect 20901 37039 21169 37047
tri 21169 37039 21177 37047 sw
rect 70802 37044 71000 37102
tri 20901 37035 20905 37039 ne
rect 20905 37036 21177 37039
rect 20905 37035 21042 37036
tri 20905 37031 20909 37035 ne
rect 20909 37031 21042 37035
tri 20909 37023 20917 37031 ne
rect 20917 37023 21042 37031
tri 20917 37015 20925 37023 ne
rect 20925 37015 21042 37023
tri 20925 37007 20933 37015 ne
rect 20933 37007 21042 37015
tri 20933 36999 20941 37007 ne
rect 20941 36999 21042 37007
tri 20941 36991 20949 36999 ne
rect 20949 36991 21042 36999
tri 20949 36983 20957 36991 ne
rect 20957 36990 21042 36991
rect 21088 37031 21177 37036
tri 21177 37031 21185 37039 sw
rect 21088 37023 21185 37031
tri 21185 37023 21193 37031 sw
rect 21088 37015 21193 37023
tri 21193 37015 21201 37023 sw
rect 21088 37007 21201 37015
tri 21201 37007 21209 37015 sw
rect 21088 36999 21209 37007
tri 21209 36999 21217 37007 sw
rect 21088 36991 21217 36999
tri 21217 36991 21225 36999 sw
rect 70802 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 21088 36990 21225 36991
rect 20957 36983 21225 36990
tri 21225 36983 21233 36991 sw
tri 20957 36975 20965 36983 ne
rect 20965 36975 21233 36983
tri 21233 36975 21241 36983 sw
tri 20965 36967 20973 36975 ne
rect 20973 36967 21241 36975
tri 21241 36967 21249 36975 sw
tri 20973 36959 20981 36967 ne
rect 20981 36959 21249 36967
tri 21249 36959 21257 36967 sw
tri 20981 36951 20989 36959 ne
rect 20989 36951 21257 36959
tri 21257 36951 21265 36959 sw
tri 20989 36943 20997 36951 ne
rect 20997 36943 21265 36951
tri 21265 36943 21273 36951 sw
tri 20997 36935 21005 36943 ne
rect 21005 36935 21273 36943
tri 21273 36935 21281 36943 sw
rect 70802 36940 71000 36998
tri 21005 36927 21013 36935 ne
rect 21013 36927 21281 36935
tri 21281 36927 21289 36935 sw
tri 21013 36919 21021 36927 ne
rect 21021 36922 21289 36927
tri 21289 36922 21294 36927 sw
rect 21021 36919 21294 36922
tri 21021 36911 21029 36919 ne
rect 21029 36914 21294 36919
tri 21294 36914 21302 36922 sw
rect 21029 36911 21302 36914
tri 21029 36908 21032 36911 ne
rect 21032 36908 21302 36911
tri 21032 36900 21040 36908 ne
rect 21040 36906 21302 36908
tri 21302 36906 21310 36914 sw
rect 21040 36904 21310 36906
rect 21040 36900 21174 36904
tri 21040 36892 21048 36900 ne
rect 21048 36892 21174 36900
tri 21048 36884 21056 36892 ne
rect 21056 36884 21174 36892
tri 21056 36876 21064 36884 ne
rect 21064 36876 21174 36884
tri 21064 36868 21072 36876 ne
rect 21072 36868 21174 36876
tri 21072 36860 21080 36868 ne
rect 21080 36860 21174 36868
tri 21080 36852 21088 36860 ne
rect 21088 36858 21174 36860
rect 21220 36898 21310 36904
tri 21310 36898 21318 36906 sw
rect 21220 36890 21318 36898
tri 21318 36890 21326 36898 sw
rect 70802 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 21220 36882 21326 36890
tri 21326 36882 21334 36890 sw
rect 21220 36874 21334 36882
tri 21334 36874 21342 36882 sw
rect 21220 36866 21342 36874
tri 21342 36866 21350 36874 sw
rect 21220 36858 21350 36866
tri 21350 36858 21358 36866 sw
rect 21088 36852 21358 36858
tri 21088 36844 21096 36852 ne
rect 21096 36850 21358 36852
tri 21358 36850 21366 36858 sw
rect 21096 36844 21366 36850
tri 21096 36836 21104 36844 ne
rect 21104 36842 21366 36844
tri 21366 36842 21374 36850 sw
rect 21104 36836 21374 36842
tri 21104 36828 21112 36836 ne
rect 21112 36834 21374 36836
tri 21374 36834 21382 36842 sw
rect 70802 36836 71000 36894
rect 21112 36828 21382 36834
tri 21112 36820 21120 36828 ne
rect 21120 36826 21382 36828
tri 21382 36826 21390 36834 sw
rect 21120 36820 21390 36826
tri 21120 36812 21128 36820 ne
rect 21128 36818 21390 36820
tri 21390 36818 21398 36826 sw
rect 21128 36812 21398 36818
tri 21128 36804 21136 36812 ne
rect 21136 36810 21398 36812
tri 21398 36810 21406 36818 sw
rect 21136 36804 21406 36810
tri 21136 36796 21144 36804 ne
rect 21144 36802 21406 36804
tri 21406 36802 21414 36810 sw
rect 21144 36796 21414 36802
tri 21144 36788 21152 36796 ne
rect 21152 36794 21414 36796
tri 21414 36794 21422 36802 sw
rect 21152 36788 21422 36794
tri 21152 36780 21160 36788 ne
rect 21160 36787 21422 36788
tri 21422 36787 21429 36794 sw
rect 70802 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21160 36780 21429 36787
tri 21160 36779 21161 36780 ne
rect 21161 36779 21429 36780
tri 21429 36779 21437 36787 sw
tri 21161 36771 21169 36779 ne
rect 21169 36772 21437 36779
rect 21169 36771 21306 36772
tri 21169 36763 21177 36771 ne
rect 21177 36763 21306 36771
tri 21177 36755 21185 36763 ne
rect 21185 36755 21306 36763
tri 21185 36747 21193 36755 ne
rect 21193 36747 21306 36755
tri 21193 36739 21201 36747 ne
rect 21201 36739 21306 36747
tri 21201 36731 21209 36739 ne
rect 21209 36731 21306 36739
tri 21209 36723 21217 36731 ne
rect 21217 36726 21306 36731
rect 21352 36771 21437 36772
tri 21437 36771 21445 36779 sw
rect 21352 36763 21445 36771
tri 21445 36763 21453 36771 sw
rect 21352 36755 21453 36763
tri 21453 36755 21461 36763 sw
rect 21352 36747 21461 36755
tri 21461 36747 21469 36755 sw
rect 21352 36739 21469 36747
tri 21469 36739 21477 36747 sw
rect 21352 36731 21477 36739
tri 21477 36731 21485 36739 sw
rect 70802 36732 71000 36790
rect 21352 36726 21485 36731
rect 21217 36723 21485 36726
tri 21485 36723 21493 36731 sw
tri 21217 36715 21225 36723 ne
rect 21225 36715 21493 36723
tri 21493 36715 21501 36723 sw
tri 21225 36707 21233 36715 ne
rect 21233 36707 21501 36715
tri 21501 36707 21509 36715 sw
tri 21233 36699 21241 36707 ne
rect 21241 36699 21509 36707
tri 21509 36699 21517 36707 sw
tri 21241 36691 21249 36699 ne
rect 21249 36691 21517 36699
tri 21517 36691 21525 36699 sw
tri 21249 36683 21257 36691 ne
rect 21257 36683 21525 36691
tri 21525 36683 21533 36691 sw
rect 70802 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
tri 21257 36675 21265 36683 ne
rect 21265 36675 21533 36683
tri 21533 36675 21541 36683 sw
tri 21265 36667 21273 36675 ne
rect 21273 36667 21541 36675
tri 21541 36667 21549 36675 sw
tri 21273 36659 21281 36667 ne
rect 21281 36659 21549 36667
tri 21549 36659 21557 36667 sw
tri 21281 36651 21289 36659 ne
rect 21289 36651 21557 36659
tri 21557 36651 21565 36659 sw
tri 21289 36650 21290 36651 ne
rect 21290 36650 21565 36651
tri 21565 36650 21566 36651 sw
tri 21290 36642 21298 36650 ne
rect 21298 36642 21566 36650
tri 21566 36642 21574 36650 sw
tri 21298 36634 21306 36642 ne
rect 21306 36640 21574 36642
rect 21306 36634 21438 36640
tri 21306 36626 21314 36634 ne
rect 21314 36626 21438 36634
tri 21314 36618 21322 36626 ne
rect 21322 36618 21438 36626
tri 21322 36610 21330 36618 ne
rect 21330 36610 21438 36618
tri 21330 36602 21338 36610 ne
rect 21338 36602 21438 36610
tri 21338 36594 21346 36602 ne
rect 21346 36594 21438 36602
rect 21484 36634 21574 36640
tri 21574 36634 21582 36642 sw
rect 21484 36626 21582 36634
tri 21582 36626 21590 36634 sw
rect 70802 36628 71000 36686
rect 21484 36618 21590 36626
tri 21590 36618 21598 36626 sw
rect 21484 36610 21598 36618
tri 21598 36610 21606 36618 sw
rect 21484 36602 21606 36610
tri 21606 36602 21614 36610 sw
rect 21484 36594 21614 36602
tri 21614 36594 21622 36602 sw
tri 21346 36586 21354 36594 ne
rect 21354 36586 21622 36594
tri 21622 36586 21630 36594 sw
tri 21354 36578 21362 36586 ne
rect 21362 36578 21630 36586
tri 21630 36578 21638 36586 sw
rect 70802 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21362 36570 21370 36578 ne
rect 21370 36570 21638 36578
tri 21638 36570 21646 36578 sw
tri 21370 36562 21378 36570 ne
rect 21378 36562 21646 36570
tri 21646 36562 21654 36570 sw
tri 21378 36554 21386 36562 ne
rect 21386 36554 21654 36562
tri 21654 36554 21662 36562 sw
tri 21386 36546 21394 36554 ne
rect 21394 36546 21662 36554
tri 21662 36546 21670 36554 sw
tri 21394 36538 21402 36546 ne
rect 21402 36538 21670 36546
tri 21670 36538 21678 36546 sw
tri 21402 36534 21406 36538 ne
rect 21406 36534 21678 36538
tri 21678 36534 21682 36538 sw
tri 21406 36530 21410 36534 ne
rect 21410 36530 21682 36534
tri 21682 36530 21686 36534 sw
tri 21410 36522 21418 36530 ne
rect 21418 36522 21686 36530
tri 21686 36522 21694 36530 sw
rect 70802 36524 71000 36582
tri 21418 36514 21426 36522 ne
rect 21426 36514 21694 36522
tri 21694 36514 21702 36522 sw
tri 21426 36506 21434 36514 ne
rect 21434 36508 21702 36514
rect 21434 36506 21570 36508
tri 21434 36498 21442 36506 ne
rect 21442 36498 21570 36506
tri 21442 36490 21450 36498 ne
rect 21450 36490 21570 36498
tri 21450 36482 21458 36490 ne
rect 21458 36482 21570 36490
tri 21458 36474 21466 36482 ne
rect 21466 36474 21570 36482
tri 21466 36466 21474 36474 ne
rect 21474 36466 21570 36474
tri 21474 36458 21482 36466 ne
rect 21482 36462 21570 36466
rect 21616 36506 21702 36508
tri 21702 36506 21710 36514 sw
rect 21616 36498 21710 36506
tri 21710 36498 21718 36506 sw
rect 21616 36490 21718 36498
tri 21718 36490 21726 36498 sw
rect 21616 36482 21726 36490
tri 21726 36482 21734 36490 sw
rect 21616 36474 21734 36482
tri 21734 36474 21742 36482 sw
rect 70802 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 21616 36466 21742 36474
tri 21742 36466 21750 36474 sw
rect 21616 36462 21750 36466
rect 21482 36458 21750 36462
tri 21750 36458 21758 36466 sw
tri 21482 36450 21490 36458 ne
rect 21490 36450 21758 36458
tri 21758 36450 21766 36458 sw
tri 21490 36442 21498 36450 ne
rect 21498 36442 21766 36450
tri 21766 36442 21774 36450 sw
tri 21498 36434 21506 36442 ne
rect 21506 36434 21774 36442
tri 21774 36434 21782 36442 sw
tri 21506 36426 21514 36434 ne
rect 21514 36426 21782 36434
tri 21782 36426 21790 36434 sw
tri 21514 36418 21522 36426 ne
rect 21522 36418 21790 36426
tri 21790 36418 21798 36426 sw
rect 70802 36420 71000 36478
tri 21522 36410 21530 36418 ne
rect 21530 36410 21798 36418
tri 21798 36410 21806 36418 sw
tri 21530 36402 21538 36410 ne
rect 21538 36409 21806 36410
tri 21806 36409 21807 36410 sw
rect 21538 36402 21807 36409
tri 21538 36401 21539 36402 ne
rect 21539 36401 21807 36402
tri 21807 36401 21815 36409 sw
tri 21539 36393 21547 36401 ne
rect 21547 36393 21815 36401
tri 21815 36393 21823 36401 sw
tri 21547 36385 21555 36393 ne
rect 21555 36385 21823 36393
tri 21823 36385 21831 36393 sw
tri 21555 36377 21563 36385 ne
rect 21563 36377 21831 36385
tri 21831 36377 21839 36385 sw
tri 21563 36369 21571 36377 ne
rect 21571 36376 21839 36377
rect 21571 36369 21702 36376
tri 21571 36361 21579 36369 ne
rect 21579 36361 21702 36369
tri 21579 36353 21587 36361 ne
rect 21587 36353 21702 36361
tri 21587 36345 21595 36353 ne
rect 21595 36345 21702 36353
tri 21595 36337 21603 36345 ne
rect 21603 36337 21702 36345
tri 21603 36329 21611 36337 ne
rect 21611 36330 21702 36337
rect 21748 36369 21839 36376
tri 21839 36369 21847 36377 sw
rect 70802 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36361 21847 36369
tri 21847 36361 21855 36369 sw
rect 21748 36353 21855 36361
tri 21855 36353 21863 36361 sw
rect 21748 36345 21863 36353
tri 21863 36345 21871 36353 sw
rect 21748 36337 21871 36345
tri 21871 36337 21879 36345 sw
rect 21748 36330 21879 36337
rect 21611 36329 21879 36330
tri 21879 36329 21887 36337 sw
tri 21611 36321 21619 36329 ne
rect 21619 36321 21887 36329
tri 21887 36321 21895 36329 sw
tri 21619 36313 21627 36321 ne
rect 21627 36313 21895 36321
tri 21895 36313 21903 36321 sw
rect 70802 36316 71000 36374
tri 21627 36305 21635 36313 ne
rect 21635 36305 21903 36313
tri 21903 36305 21911 36313 sw
tri 21635 36297 21643 36305 ne
rect 21643 36297 21911 36305
tri 21911 36297 21919 36305 sw
tri 21643 36289 21651 36297 ne
rect 21651 36289 21919 36297
tri 21919 36289 21927 36297 sw
tri 21651 36281 21659 36289 ne
rect 21659 36281 21927 36289
tri 21927 36281 21935 36289 sw
tri 21659 36273 21667 36281 ne
rect 21667 36273 21935 36281
tri 21935 36273 21943 36281 sw
tri 21667 36267 21673 36273 ne
rect 21673 36267 21943 36273
tri 21943 36267 21949 36273 sw
rect 70802 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
tri 21673 36259 21681 36267 ne
rect 21681 36259 21949 36267
tri 21949 36259 21957 36267 sw
tri 21681 36254 21686 36259 ne
rect 21686 36254 21957 36259
tri 21686 36251 21689 36254 ne
rect 21689 36251 21957 36254
tri 21957 36251 21965 36259 sw
tri 21689 36243 21697 36251 ne
rect 21697 36244 21965 36251
rect 21697 36243 21834 36244
tri 21697 36235 21705 36243 ne
rect 21705 36235 21834 36243
tri 21705 36227 21713 36235 ne
rect 21713 36227 21834 36235
tri 21713 36219 21721 36227 ne
rect 21721 36219 21834 36227
tri 21721 36211 21729 36219 ne
rect 21729 36211 21834 36219
tri 21729 36203 21737 36211 ne
rect 21737 36203 21834 36211
tri 21737 36195 21745 36203 ne
rect 21745 36198 21834 36203
rect 21880 36243 21965 36244
tri 21965 36243 21973 36251 sw
rect 21880 36235 21973 36243
tri 21973 36235 21981 36243 sw
rect 21880 36227 21981 36235
tri 21981 36227 21989 36235 sw
rect 21880 36219 21989 36227
tri 21989 36219 21997 36227 sw
rect 21880 36211 21997 36219
tri 21997 36211 22005 36219 sw
rect 70802 36212 71000 36270
rect 21880 36203 22005 36211
tri 22005 36203 22013 36211 sw
rect 21880 36198 22013 36203
rect 21745 36195 22013 36198
tri 22013 36195 22021 36203 sw
tri 21745 36187 21753 36195 ne
rect 21753 36187 22021 36195
tri 22021 36187 22029 36195 sw
tri 21753 36179 21761 36187 ne
rect 21761 36179 22029 36187
tri 22029 36179 22037 36187 sw
tri 21761 36171 21769 36179 ne
rect 21769 36171 22037 36179
tri 22037 36171 22045 36179 sw
tri 21769 36163 21777 36171 ne
rect 21777 36163 22045 36171
tri 22045 36163 22053 36171 sw
rect 70802 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21777 36155 21785 36163 ne
rect 21785 36155 22053 36163
tri 22053 36155 22061 36163 sw
tri 21785 36147 21793 36155 ne
rect 21793 36147 22061 36155
tri 22061 36147 22069 36155 sw
tri 21793 36139 21801 36147 ne
rect 21801 36139 22069 36147
tri 22069 36139 22077 36147 sw
tri 21801 36131 21809 36139 ne
rect 21809 36131 22077 36139
tri 22077 36131 22085 36139 sw
tri 21809 36123 21817 36131 ne
rect 21817 36123 22085 36131
tri 22085 36123 22093 36131 sw
tri 21817 36115 21825 36123 ne
rect 21825 36115 22093 36123
tri 22093 36115 22101 36123 sw
tri 21825 36107 21833 36115 ne
rect 21833 36112 22101 36115
rect 21833 36107 21966 36112
tri 21833 36099 21841 36107 ne
rect 21841 36099 21966 36107
tri 21841 36091 21849 36099 ne
rect 21849 36091 21966 36099
tri 21849 36083 21857 36091 ne
rect 21857 36083 21966 36091
tri 21857 36075 21865 36083 ne
rect 21865 36075 21966 36083
tri 21865 36067 21873 36075 ne
rect 21873 36067 21966 36075
tri 21873 36059 21881 36067 ne
rect 21881 36066 21966 36067
rect 22012 36107 22101 36112
tri 22101 36107 22109 36115 sw
rect 70802 36108 71000 36166
rect 22012 36099 22109 36107
tri 22109 36099 22117 36107 sw
rect 22012 36091 22117 36099
tri 22117 36091 22125 36099 sw
rect 22012 36083 22125 36091
tri 22125 36083 22133 36091 sw
rect 22012 36075 22133 36083
tri 22133 36075 22141 36083 sw
rect 22012 36067 22141 36075
tri 22141 36067 22149 36075 sw
rect 22012 36066 22149 36067
rect 21881 36065 22149 36066
tri 22149 36065 22151 36067 sw
rect 21881 36059 22151 36065
tri 21881 36054 21886 36059 ne
rect 21886 36057 22151 36059
tri 22151 36057 22159 36065 sw
rect 70802 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
rect 21886 36054 22159 36057
tri 21886 36046 21894 36054 ne
rect 21894 36049 22159 36054
tri 22159 36049 22167 36057 sw
rect 21894 36046 22167 36049
tri 21894 36038 21902 36046 ne
rect 21902 36041 22167 36046
tri 22167 36041 22175 36049 sw
rect 21902 36038 22175 36041
tri 21902 36030 21910 36038 ne
rect 21910 36033 22175 36038
tri 22175 36033 22183 36041 sw
rect 21910 36030 22183 36033
tri 21910 36022 21918 36030 ne
rect 21918 36025 22183 36030
tri 22183 36025 22191 36033 sw
rect 21918 36022 22191 36025
tri 21918 36014 21926 36022 ne
rect 21926 36017 22191 36022
tri 22191 36017 22199 36025 sw
rect 21926 36014 22199 36017
tri 21926 36006 21934 36014 ne
rect 21934 36009 22199 36014
tri 22199 36009 22207 36017 sw
rect 21934 36006 22207 36009
tri 21934 35998 21942 36006 ne
rect 21942 36001 22207 36006
tri 22207 36001 22215 36009 sw
rect 70802 36004 71000 36062
rect 21942 35998 22215 36001
tri 21942 35990 21950 35998 ne
rect 21950 35993 22215 35998
tri 22215 35993 22223 36001 sw
rect 21950 35990 22223 35993
tri 21950 35982 21958 35990 ne
rect 21958 35985 22223 35990
tri 22223 35985 22231 35993 sw
rect 21958 35982 22231 35985
tri 21958 35974 21966 35982 ne
rect 21966 35980 22231 35982
rect 21966 35974 22098 35980
tri 21966 35966 21974 35974 ne
rect 21974 35966 22098 35974
tri 21974 35958 21982 35966 ne
rect 21982 35958 22098 35966
tri 21982 35950 21990 35958 ne
rect 21990 35950 22098 35958
tri 21990 35942 21998 35950 ne
rect 21998 35942 22098 35950
tri 21998 35934 22006 35942 ne
rect 22006 35934 22098 35942
rect 22144 35977 22231 35980
tri 22231 35977 22239 35985 sw
rect 22144 35969 22239 35977
tri 22239 35969 22247 35977 sw
rect 22144 35961 22247 35969
tri 22247 35961 22255 35969 sw
rect 22144 35953 22255 35961
tri 22255 35953 22263 35961 sw
rect 70802 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22144 35948 22263 35953
tri 22263 35948 22268 35953 sw
rect 22144 35940 22268 35948
tri 22268 35940 22276 35948 sw
rect 22144 35934 22276 35940
tri 22006 35926 22014 35934 ne
rect 22014 35932 22276 35934
tri 22276 35932 22284 35940 sw
rect 22014 35926 22284 35932
tri 22014 35918 22022 35926 ne
rect 22022 35924 22284 35926
tri 22284 35924 22292 35932 sw
rect 22022 35918 22292 35924
tri 22022 35915 22025 35918 ne
rect 22025 35916 22292 35918
tri 22292 35916 22300 35924 sw
rect 22025 35915 22300 35916
tri 22025 35907 22033 35915 ne
rect 22033 35908 22300 35915
tri 22300 35908 22308 35916 sw
rect 22033 35907 22308 35908
tri 22033 35899 22041 35907 ne
rect 22041 35900 22308 35907
tri 22308 35900 22316 35908 sw
rect 70802 35900 71000 35958
rect 22041 35899 22316 35900
tri 22041 35891 22049 35899 ne
rect 22049 35892 22316 35899
tri 22316 35892 22324 35900 sw
rect 22049 35891 22324 35892
tri 22049 35883 22057 35891 ne
rect 22057 35884 22324 35891
tri 22324 35884 22332 35892 sw
rect 22057 35883 22332 35884
tri 22057 35875 22065 35883 ne
rect 22065 35876 22332 35883
tri 22332 35876 22340 35884 sw
rect 22065 35875 22340 35876
tri 22065 35867 22073 35875 ne
rect 22073 35868 22340 35875
tri 22340 35868 22348 35876 sw
rect 22073 35867 22348 35868
tri 22073 35859 22081 35867 ne
rect 22081 35860 22348 35867
tri 22348 35860 22356 35868 sw
rect 22081 35859 22356 35860
tri 22081 35851 22089 35859 ne
rect 22089 35852 22356 35859
tri 22356 35852 22364 35860 sw
rect 70802 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 22089 35851 22364 35852
tri 22089 35843 22097 35851 ne
rect 22097 35848 22364 35851
rect 22097 35843 22230 35848
tri 22097 35835 22105 35843 ne
rect 22105 35835 22230 35843
tri 22105 35827 22113 35835 ne
rect 22113 35827 22230 35835
tri 22113 35819 22121 35827 ne
rect 22121 35819 22230 35827
tri 22121 35811 22129 35819 ne
rect 22129 35811 22230 35819
tri 22129 35803 22137 35811 ne
rect 22137 35803 22230 35811
tri 22137 35795 22145 35803 ne
rect 22145 35802 22230 35803
rect 22276 35844 22364 35848
tri 22364 35844 22372 35852 sw
rect 22276 35836 22372 35844
tri 22372 35836 22380 35844 sw
rect 22276 35828 22380 35836
tri 22380 35828 22388 35836 sw
rect 22276 35820 22388 35828
tri 22388 35820 22396 35828 sw
rect 22276 35812 22396 35820
tri 22396 35812 22404 35820 sw
rect 22276 35811 22404 35812
tri 22404 35811 22405 35812 sw
rect 22276 35803 22405 35811
tri 22405 35803 22413 35811 sw
rect 22276 35802 22413 35803
rect 22145 35795 22413 35802
tri 22413 35795 22421 35803 sw
rect 70802 35796 71000 35854
tri 22145 35789 22151 35795 ne
rect 22151 35789 22421 35795
tri 22151 35781 22159 35789 ne
rect 22159 35787 22421 35789
tri 22421 35787 22429 35795 sw
rect 22159 35781 22429 35787
tri 22159 35773 22167 35781 ne
rect 22167 35779 22429 35781
tri 22429 35779 22437 35787 sw
rect 22167 35773 22437 35779
tri 22167 35765 22175 35773 ne
rect 22175 35771 22437 35773
tri 22437 35771 22445 35779 sw
rect 22175 35765 22445 35771
tri 22175 35757 22183 35765 ne
rect 22183 35763 22445 35765
tri 22445 35763 22453 35771 sw
rect 22183 35757 22453 35763
tri 22183 35749 22191 35757 ne
rect 22191 35755 22453 35757
tri 22453 35755 22461 35763 sw
rect 22191 35749 22461 35755
tri 22191 35741 22199 35749 ne
rect 22199 35747 22461 35749
tri 22461 35747 22469 35755 sw
rect 70802 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
rect 22199 35741 22469 35747
tri 22199 35733 22207 35741 ne
rect 22207 35739 22469 35741
tri 22469 35739 22477 35747 sw
rect 22207 35733 22477 35739
tri 22207 35725 22215 35733 ne
rect 22215 35731 22477 35733
tri 22477 35731 22485 35739 sw
rect 22215 35729 22485 35731
tri 22485 35729 22487 35731 sw
rect 22215 35725 22487 35729
tri 22215 35717 22223 35725 ne
rect 22223 35723 22487 35725
tri 22487 35723 22493 35729 sw
rect 22223 35717 22493 35723
tri 22223 35709 22231 35717 ne
rect 22231 35716 22493 35717
rect 22231 35709 22362 35716
tri 22231 35701 22239 35709 ne
rect 22239 35701 22362 35709
tri 22239 35693 22247 35701 ne
rect 22247 35693 22362 35701
tri 22247 35685 22255 35693 ne
rect 22255 35685 22362 35693
tri 22255 35677 22263 35685 ne
rect 22263 35677 22362 35685
tri 22263 35669 22271 35677 ne
rect 22271 35670 22362 35677
rect 22408 35715 22493 35716
tri 22493 35715 22501 35723 sw
rect 22408 35707 22501 35715
tri 22501 35707 22509 35715 sw
rect 22408 35699 22509 35707
tri 22509 35699 22517 35707 sw
rect 22408 35691 22517 35699
tri 22517 35691 22525 35699 sw
rect 70802 35692 71000 35750
rect 22408 35683 22525 35691
tri 22525 35683 22533 35691 sw
rect 22408 35675 22533 35683
tri 22533 35675 22541 35683 sw
rect 22408 35670 22541 35675
rect 22271 35669 22541 35670
tri 22271 35661 22279 35669 ne
rect 22279 35667 22541 35669
tri 22541 35667 22549 35675 sw
rect 22279 35661 22549 35667
tri 22279 35653 22287 35661 ne
rect 22287 35659 22549 35661
tri 22549 35659 22557 35667 sw
rect 22287 35653 22557 35659
tri 22287 35645 22295 35653 ne
rect 22295 35651 22557 35653
tri 22557 35651 22565 35659 sw
rect 22295 35645 22565 35651
tri 22295 35637 22303 35645 ne
rect 22303 35643 22565 35645
tri 22565 35643 22573 35651 sw
rect 70802 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 22303 35637 22573 35643
tri 22303 35629 22311 35637 ne
rect 22311 35635 22573 35637
tri 22573 35635 22581 35643 sw
rect 22311 35629 22581 35635
tri 22311 35621 22319 35629 ne
rect 22319 35627 22581 35629
tri 22581 35627 22589 35635 sw
rect 22319 35621 22589 35627
tri 22319 35613 22327 35621 ne
rect 22327 35619 22589 35621
tri 22589 35619 22597 35627 sw
rect 22327 35613 22597 35619
tri 22327 35605 22335 35613 ne
rect 22335 35611 22597 35613
tri 22597 35611 22605 35619 sw
rect 22335 35605 22605 35611
tri 22335 35597 22343 35605 ne
rect 22343 35603 22605 35605
tri 22605 35603 22613 35611 sw
rect 22343 35597 22613 35603
tri 22343 35589 22351 35597 ne
rect 22351 35595 22613 35597
tri 22613 35595 22621 35603 sw
rect 22351 35593 22621 35595
tri 22621 35593 22623 35595 sw
rect 22351 35589 22623 35593
tri 22351 35581 22359 35589 ne
rect 22359 35585 22623 35589
tri 22623 35585 22631 35593 sw
rect 70802 35588 71000 35646
rect 22359 35584 22631 35585
rect 22359 35581 22494 35584
tri 22359 35573 22367 35581 ne
rect 22367 35573 22494 35581
tri 22367 35565 22375 35573 ne
rect 22375 35565 22494 35573
tri 22375 35557 22383 35565 ne
rect 22383 35557 22494 35565
tri 22383 35549 22391 35557 ne
rect 22391 35549 22494 35557
tri 22391 35541 22399 35549 ne
rect 22399 35541 22494 35549
tri 22399 35537 22403 35541 ne
rect 22403 35538 22494 35541
rect 22540 35577 22631 35584
tri 22631 35577 22639 35585 sw
rect 22540 35569 22639 35577
tri 22639 35569 22647 35577 sw
rect 22540 35561 22647 35569
tri 22647 35561 22655 35569 sw
rect 22540 35553 22655 35561
tri 22655 35553 22663 35561 sw
rect 22540 35545 22663 35553
tri 22663 35545 22671 35553 sw
rect 22540 35538 22671 35545
rect 22403 35537 22671 35538
tri 22671 35537 22679 35545 sw
rect 70802 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
tri 22403 35529 22411 35537 ne
rect 22411 35529 22679 35537
tri 22679 35529 22687 35537 sw
tri 22411 35521 22419 35529 ne
rect 22419 35521 22687 35529
tri 22687 35521 22695 35529 sw
tri 22419 35513 22427 35521 ne
rect 22427 35513 22695 35521
tri 22695 35513 22703 35521 sw
tri 22427 35505 22435 35513 ne
rect 22435 35505 22703 35513
tri 22703 35505 22711 35513 sw
tri 22435 35497 22443 35505 ne
rect 22443 35497 22711 35505
tri 22711 35497 22719 35505 sw
tri 22443 35489 22451 35497 ne
rect 22451 35489 22719 35497
tri 22719 35489 22727 35497 sw
tri 22451 35481 22459 35489 ne
rect 22459 35481 22727 35489
tri 22727 35481 22735 35489 sw
rect 70802 35484 71000 35542
tri 22459 35473 22467 35481 ne
rect 22467 35473 22735 35481
tri 22735 35473 22743 35481 sw
tri 22467 35465 22475 35473 ne
rect 22475 35465 22743 35473
tri 22743 35465 22751 35473 sw
tri 22475 35457 22483 35465 ne
rect 22483 35457 22751 35465
tri 22751 35457 22759 35465 sw
tri 22483 35453 22487 35457 ne
rect 22487 35453 22759 35457
tri 22759 35453 22763 35457 sw
tri 22487 35449 22491 35453 ne
rect 22491 35452 22763 35453
rect 22491 35449 22626 35452
tri 22491 35441 22499 35449 ne
rect 22499 35441 22626 35449
tri 22499 35433 22507 35441 ne
rect 22507 35433 22626 35441
tri 22507 35425 22515 35433 ne
rect 22515 35425 22626 35433
tri 22515 35417 22523 35425 ne
rect 22523 35417 22626 35425
tri 22523 35409 22531 35417 ne
rect 22531 35409 22626 35417
tri 22531 35401 22539 35409 ne
rect 22539 35406 22626 35409
rect 22672 35449 22763 35452
tri 22763 35449 22767 35453 sw
rect 22672 35441 22767 35449
tri 22767 35441 22775 35449 sw
rect 22672 35433 22775 35441
tri 22775 35433 22783 35441 sw
rect 70802 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35425 22783 35433
tri 22783 35425 22791 35433 sw
rect 22672 35417 22791 35425
tri 22791 35417 22799 35425 sw
rect 22672 35409 22799 35417
tri 22799 35409 22807 35417 sw
rect 22672 35406 22807 35409
rect 22539 35401 22807 35406
tri 22807 35401 22815 35409 sw
tri 22539 35393 22547 35401 ne
rect 22547 35393 22815 35401
tri 22815 35393 22823 35401 sw
tri 22547 35385 22555 35393 ne
rect 22555 35385 22823 35393
tri 22823 35385 22831 35393 sw
tri 22555 35377 22563 35385 ne
rect 22563 35377 22831 35385
tri 22831 35377 22839 35385 sw
rect 70802 35380 71000 35438
tri 22563 35369 22571 35377 ne
rect 22571 35369 22839 35377
tri 22839 35369 22847 35377 sw
tri 22571 35361 22579 35369 ne
rect 22579 35361 22847 35369
tri 22847 35361 22855 35369 sw
tri 22579 35353 22587 35361 ne
rect 22587 35353 22855 35361
tri 22855 35353 22863 35361 sw
tri 22587 35345 22595 35353 ne
rect 22595 35345 22863 35353
tri 22863 35345 22871 35353 sw
tri 22595 35337 22603 35345 ne
rect 22603 35337 22871 35345
tri 22871 35337 22879 35345 sw
tri 22603 35329 22611 35337 ne
rect 22611 35334 22879 35337
tri 22879 35334 22882 35337 sw
rect 70802 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22611 35329 22882 35334
tri 22611 35321 22619 35329 ne
rect 22619 35326 22882 35329
tri 22882 35326 22890 35334 sw
rect 22619 35321 22890 35326
tri 22619 35314 22626 35321 ne
rect 22626 35320 22890 35321
rect 22626 35314 22758 35320
tri 22626 35306 22634 35314 ne
rect 22634 35306 22758 35314
tri 22634 35298 22642 35306 ne
rect 22642 35298 22758 35306
tri 22642 35290 22650 35298 ne
rect 22650 35290 22758 35298
tri 22650 35282 22658 35290 ne
rect 22658 35282 22758 35290
tri 22658 35274 22666 35282 ne
rect 22666 35274 22758 35282
rect 22804 35318 22890 35320
tri 22890 35318 22898 35326 sw
rect 22804 35310 22898 35318
tri 22898 35310 22906 35318 sw
rect 22804 35302 22906 35310
tri 22906 35302 22914 35310 sw
rect 22804 35294 22914 35302
tri 22914 35294 22922 35302 sw
rect 22804 35286 22922 35294
tri 22922 35286 22930 35294 sw
rect 22804 35278 22930 35286
tri 22930 35278 22938 35286 sw
rect 22804 35274 22938 35278
tri 22666 35266 22674 35274 ne
rect 22674 35270 22938 35274
tri 22938 35270 22946 35278 sw
rect 70802 35276 71000 35334
rect 22674 35266 22946 35270
tri 22674 35258 22682 35266 ne
rect 22682 35262 22946 35266
tri 22946 35262 22954 35270 sw
rect 22682 35258 22954 35262
tri 22682 35250 22690 35258 ne
rect 22690 35254 22954 35258
tri 22954 35254 22962 35262 sw
rect 22690 35250 22962 35254
tri 22690 35242 22698 35250 ne
rect 22698 35246 22962 35250
tri 22962 35246 22970 35254 sw
rect 22698 35242 22970 35246
tri 22698 35234 22706 35242 ne
rect 22706 35238 22970 35242
tri 22970 35238 22978 35246 sw
rect 22706 35234 22978 35238
tri 22706 35226 22714 35234 ne
rect 22714 35230 22978 35234
tri 22978 35230 22986 35238 sw
rect 70802 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
rect 22714 35226 22986 35230
tri 22714 35218 22722 35226 ne
rect 22722 35222 22986 35226
tri 22986 35222 22994 35230 sw
rect 22722 35218 22994 35222
tri 22722 35210 22730 35218 ne
rect 22730 35214 22994 35218
tri 22994 35214 23002 35222 sw
rect 22730 35210 23002 35214
tri 22730 35202 22738 35210 ne
rect 22738 35207 23002 35210
tri 23002 35207 23009 35214 sw
rect 22738 35202 23009 35207
tri 22738 35194 22746 35202 ne
rect 22746 35199 23009 35202
tri 23009 35199 23017 35207 sw
rect 22746 35194 23017 35199
tri 22746 35186 22754 35194 ne
rect 22754 35191 23017 35194
tri 23017 35191 23025 35199 sw
rect 22754 35188 23025 35191
rect 22754 35186 22890 35188
tri 22754 35182 22758 35186 ne
rect 22758 35182 22890 35186
tri 22758 35178 22762 35182 ne
rect 22762 35178 22890 35182
tri 22762 35170 22770 35178 ne
rect 22770 35170 22890 35178
tri 22770 35162 22778 35170 ne
rect 22778 35162 22890 35170
tri 22778 35154 22786 35162 ne
rect 22786 35154 22890 35162
tri 22786 35146 22794 35154 ne
rect 22794 35146 22890 35154
tri 22794 35138 22802 35146 ne
rect 22802 35142 22890 35146
rect 22936 35183 23025 35188
tri 23025 35183 23033 35191 sw
rect 22936 35178 23033 35183
tri 23033 35178 23038 35183 sw
rect 22936 35170 23038 35178
tri 23038 35170 23046 35178 sw
rect 70802 35172 71000 35230
rect 22936 35162 23046 35170
tri 23046 35162 23054 35170 sw
rect 22936 35154 23054 35162
tri 23054 35154 23062 35162 sw
rect 22936 35146 23062 35154
tri 23062 35146 23070 35154 sw
rect 22936 35142 23070 35146
rect 22802 35138 23070 35142
tri 23070 35138 23078 35146 sw
tri 22802 35130 22810 35138 ne
rect 22810 35130 23078 35138
tri 23078 35130 23086 35138 sw
tri 22810 35122 22818 35130 ne
rect 22818 35126 23086 35130
tri 23086 35126 23090 35130 sw
rect 70802 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
rect 22818 35122 23090 35126
tri 22818 35118 22822 35122 ne
rect 22822 35118 23090 35122
tri 23090 35118 23098 35126 sw
tri 22822 35110 22830 35118 ne
rect 22830 35110 23098 35118
tri 23098 35110 23106 35118 sw
tri 22830 35102 22838 35110 ne
rect 22838 35102 23106 35110
tri 23106 35102 23114 35110 sw
tri 22838 35094 22846 35102 ne
rect 22846 35094 23114 35102
tri 23114 35094 23122 35102 sw
tri 22846 35086 22854 35094 ne
rect 22854 35086 23122 35094
tri 23122 35086 23130 35094 sw
tri 22854 35078 22862 35086 ne
rect 22862 35078 23130 35086
tri 23130 35078 23138 35086 sw
tri 22862 35070 22870 35078 ne
rect 22870 35070 23138 35078
tri 23138 35070 23146 35078 sw
tri 22870 35062 22878 35070 ne
rect 22878 35062 23146 35070
tri 23146 35062 23154 35070 sw
rect 70802 35068 71000 35126
tri 22878 35054 22886 35062 ne
rect 22886 35056 23154 35062
rect 22886 35054 23022 35056
tri 22886 35046 22894 35054 ne
rect 22894 35046 23022 35054
tri 22894 35038 22902 35046 ne
rect 22902 35038 23022 35046
tri 22902 35030 22910 35038 ne
rect 22910 35030 23022 35038
tri 22910 35022 22918 35030 ne
rect 22918 35022 23022 35030
tri 22918 35014 22926 35022 ne
rect 22926 35014 23022 35022
tri 22926 35006 22934 35014 ne
rect 22934 35010 23022 35014
rect 23068 35054 23154 35056
tri 23154 35054 23162 35062 sw
rect 23068 35046 23162 35054
tri 23162 35046 23170 35054 sw
rect 23068 35038 23170 35046
tri 23170 35038 23178 35046 sw
rect 23068 35030 23178 35038
tri 23178 35030 23186 35038 sw
rect 23068 35022 23186 35030
tri 23186 35022 23194 35030 sw
rect 70802 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 23068 35014 23194 35022
tri 23194 35014 23202 35022 sw
rect 23068 35010 23202 35014
tri 23202 35010 23206 35014 sw
rect 22934 35006 23206 35010
tri 22934 34998 22942 35006 ne
rect 22942 35002 23206 35006
tri 23206 35002 23214 35010 sw
rect 22942 34998 23214 35002
tri 22942 34990 22950 34998 ne
rect 22950 34994 23214 34998
tri 23214 34994 23222 35002 sw
rect 22950 34990 23222 34994
tri 22950 34987 22953 34990 ne
rect 22953 34987 23222 34990
tri 22953 34979 22961 34987 ne
rect 22961 34986 23222 34987
tri 23222 34986 23230 34994 sw
rect 22961 34979 23230 34986
tri 22961 34971 22969 34979 ne
rect 22969 34978 23230 34979
tri 23230 34978 23238 34986 sw
rect 22969 34971 23238 34978
tri 22969 34963 22977 34971 ne
rect 22977 34970 23238 34971
tri 23238 34970 23246 34978 sw
rect 22977 34963 23246 34970
tri 22977 34955 22985 34963 ne
rect 22985 34962 23246 34963
tri 23246 34962 23254 34970 sw
rect 70802 34964 71000 35022
rect 22985 34955 23254 34962
tri 22985 34947 22993 34955 ne
rect 22993 34954 23254 34955
tri 23254 34954 23262 34962 sw
rect 22993 34947 23262 34954
tri 22993 34939 23001 34947 ne
rect 23001 34946 23262 34947
tri 23262 34946 23270 34954 sw
rect 23001 34939 23270 34946
tri 23001 34931 23009 34939 ne
rect 23009 34938 23270 34939
tri 23270 34938 23278 34946 sw
rect 23009 34931 23278 34938
tri 23009 34923 23017 34931 ne
rect 23017 34930 23278 34931
tri 23278 34930 23286 34938 sw
rect 23017 34924 23286 34930
rect 23017 34923 23154 34924
tri 23017 34915 23025 34923 ne
rect 23025 34915 23154 34923
tri 23025 34907 23033 34915 ne
rect 23033 34907 23154 34915
tri 23033 34899 23041 34907 ne
rect 23041 34899 23154 34907
tri 23041 34891 23049 34899 ne
rect 23049 34891 23154 34899
tri 23049 34883 23057 34891 ne
rect 23057 34883 23154 34891
tri 23057 34875 23065 34883 ne
rect 23065 34878 23154 34883
rect 23200 34923 23286 34924
tri 23286 34923 23293 34930 sw
rect 23200 34915 23293 34923
tri 23293 34915 23301 34923 sw
rect 70802 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34907 23301 34915
tri 23301 34907 23309 34915 sw
rect 23200 34899 23309 34907
tri 23309 34899 23317 34907 sw
rect 23200 34891 23317 34899
tri 23317 34891 23325 34899 sw
rect 23200 34883 23325 34891
tri 23325 34883 23333 34891 sw
rect 23200 34878 23333 34883
rect 23065 34875 23333 34878
tri 23333 34875 23341 34883 sw
tri 23065 34867 23073 34875 ne
rect 23073 34867 23341 34875
tri 23341 34867 23349 34875 sw
tri 23073 34859 23081 34867 ne
rect 23081 34859 23349 34867
tri 23349 34859 23357 34867 sw
rect 70802 34860 71000 34918
tri 23081 34851 23089 34859 ne
rect 23089 34851 23357 34859
tri 23357 34851 23365 34859 sw
tri 23089 34849 23091 34851 ne
rect 23091 34849 23365 34851
tri 23091 34841 23099 34849 ne
rect 23099 34843 23365 34849
tri 23365 34843 23373 34851 sw
rect 23099 34841 23373 34843
tri 23099 34833 23107 34841 ne
rect 23107 34835 23373 34841
tri 23373 34835 23381 34843 sw
rect 23107 34833 23381 34835
tri 23107 34825 23115 34833 ne
rect 23115 34827 23381 34833
tri 23381 34827 23389 34835 sw
rect 23115 34825 23389 34827
tri 23115 34817 23123 34825 ne
rect 23123 34819 23389 34825
tri 23389 34819 23397 34827 sw
rect 23123 34817 23397 34819
tri 23123 34809 23131 34817 ne
rect 23131 34811 23397 34817
tri 23397 34811 23405 34819 sw
rect 70802 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23131 34809 23405 34811
tri 23131 34801 23139 34809 ne
rect 23139 34803 23405 34809
tri 23405 34803 23413 34811 sw
rect 23139 34801 23413 34803
tri 23139 34793 23147 34801 ne
rect 23147 34800 23413 34801
tri 23413 34800 23416 34803 sw
rect 23147 34793 23416 34800
tri 23147 34785 23155 34793 ne
rect 23155 34792 23416 34793
tri 23416 34792 23424 34800 sw
rect 23155 34785 23286 34792
tri 23155 34777 23163 34785 ne
rect 23163 34777 23286 34785
tri 23163 34769 23171 34777 ne
rect 23171 34769 23286 34777
tri 23171 34761 23179 34769 ne
rect 23179 34761 23286 34769
tri 23179 34753 23187 34761 ne
rect 23187 34753 23286 34761
tri 23187 34745 23195 34753 ne
rect 23195 34746 23286 34753
rect 23332 34784 23424 34792
tri 23424 34784 23432 34792 sw
rect 23332 34776 23432 34784
tri 23432 34776 23440 34784 sw
rect 23332 34768 23440 34776
tri 23440 34768 23448 34776 sw
rect 23332 34760 23448 34768
tri 23448 34760 23456 34768 sw
rect 23332 34752 23456 34760
tri 23456 34752 23464 34760 sw
rect 70802 34756 71000 34814
rect 23332 34746 23464 34752
rect 23195 34745 23464 34746
tri 23195 34737 23203 34745 ne
rect 23203 34744 23464 34745
tri 23464 34744 23472 34752 sw
rect 23203 34737 23472 34744
tri 23203 34730 23210 34737 ne
rect 23210 34736 23472 34737
tri 23472 34736 23480 34744 sw
rect 23210 34730 23480 34736
tri 23210 34722 23218 34730 ne
rect 23218 34728 23480 34730
tri 23480 34728 23488 34736 sw
rect 23218 34722 23488 34728
tri 23218 34714 23226 34722 ne
rect 23226 34720 23488 34722
tri 23488 34720 23496 34728 sw
rect 23226 34714 23496 34720
tri 23226 34706 23234 34714 ne
rect 23234 34712 23496 34714
tri 23496 34712 23504 34720 sw
rect 23234 34706 23504 34712
tri 23234 34698 23242 34706 ne
rect 23242 34704 23504 34706
tri 23504 34704 23512 34712 sw
rect 70802 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
rect 23242 34698 23512 34704
tri 23242 34690 23250 34698 ne
rect 23250 34696 23512 34698
tri 23512 34696 23520 34704 sw
rect 23250 34690 23520 34696
tri 23250 34682 23258 34690 ne
rect 23258 34688 23520 34690
tri 23520 34688 23528 34696 sw
rect 23258 34687 23528 34688
tri 23528 34687 23529 34688 sw
rect 23258 34682 23529 34687
tri 23258 34674 23266 34682 ne
rect 23266 34679 23529 34682
tri 23529 34679 23537 34687 sw
rect 23266 34674 23537 34679
tri 23266 34670 23270 34674 ne
rect 23270 34671 23537 34674
tri 23537 34671 23545 34679 sw
rect 23270 34670 23545 34671
tri 23270 34666 23274 34670 ne
rect 23274 34666 23545 34670
tri 23545 34666 23550 34671 sw
tri 23274 34658 23282 34666 ne
rect 23282 34663 23550 34666
tri 23550 34663 23553 34666 sw
rect 23282 34660 23553 34663
rect 23282 34658 23418 34660
tri 23282 34650 23290 34658 ne
rect 23290 34650 23418 34658
tri 23290 34642 23298 34650 ne
rect 23298 34642 23418 34650
tri 23298 34634 23306 34642 ne
rect 23306 34634 23418 34642
tri 23306 34626 23314 34634 ne
rect 23314 34626 23418 34634
tri 23314 34618 23322 34626 ne
rect 23322 34618 23418 34626
tri 23322 34610 23330 34618 ne
rect 23330 34614 23418 34618
rect 23464 34655 23553 34660
tri 23553 34655 23561 34663 sw
rect 23464 34647 23561 34655
tri 23561 34647 23569 34655 sw
rect 70802 34652 71000 34710
rect 23464 34639 23569 34647
tri 23569 34639 23577 34647 sw
rect 23464 34631 23577 34639
tri 23577 34631 23585 34639 sw
rect 23464 34623 23585 34631
tri 23585 34623 23593 34631 sw
rect 23464 34617 23593 34623
tri 23593 34617 23599 34623 sw
rect 23464 34614 23599 34617
rect 23330 34610 23599 34614
tri 23330 34602 23338 34610 ne
rect 23338 34609 23599 34610
tri 23599 34609 23607 34617 sw
rect 23338 34602 23607 34609
tri 23338 34594 23346 34602 ne
rect 23346 34601 23607 34602
tri 23607 34601 23615 34609 sw
rect 70802 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 23346 34594 23615 34601
tri 23346 34590 23350 34594 ne
rect 23350 34593 23615 34594
tri 23615 34593 23623 34601 sw
rect 23350 34590 23623 34593
tri 23350 34582 23358 34590 ne
rect 23358 34585 23623 34590
tri 23623 34585 23631 34593 sw
rect 23358 34582 23631 34585
tri 23358 34574 23366 34582 ne
rect 23366 34577 23631 34582
tri 23631 34577 23639 34585 sw
rect 23366 34574 23639 34577
tri 23366 34566 23374 34574 ne
rect 23374 34569 23639 34574
tri 23639 34569 23647 34577 sw
rect 23374 34566 23647 34569
tri 23374 34558 23382 34566 ne
rect 23382 34561 23647 34566
tri 23647 34561 23655 34569 sw
rect 23382 34558 23655 34561
tri 23382 34550 23390 34558 ne
rect 23390 34553 23655 34558
tri 23655 34553 23663 34561 sw
rect 23390 34550 23663 34553
tri 23390 34542 23398 34550 ne
rect 23398 34545 23663 34550
tri 23663 34545 23671 34553 sw
rect 70802 34548 71000 34606
rect 23398 34542 23671 34545
tri 23398 34534 23406 34542 ne
rect 23406 34537 23671 34542
tri 23671 34537 23679 34545 sw
rect 23406 34534 23679 34537
tri 23406 34526 23414 34534 ne
rect 23414 34529 23679 34534
tri 23679 34529 23687 34537 sw
rect 23414 34528 23687 34529
rect 23414 34526 23550 34528
tri 23414 34518 23422 34526 ne
rect 23422 34518 23550 34526
tri 23422 34510 23430 34518 ne
rect 23430 34510 23550 34518
tri 23430 34502 23438 34510 ne
rect 23438 34502 23550 34510
tri 23438 34494 23446 34502 ne
rect 23446 34494 23550 34502
tri 23446 34486 23454 34494 ne
rect 23454 34486 23550 34494
tri 23454 34478 23462 34486 ne
rect 23462 34482 23550 34486
rect 23596 34521 23687 34528
tri 23687 34521 23695 34529 sw
rect 23596 34513 23695 34521
tri 23695 34513 23703 34521 sw
rect 23596 34505 23703 34513
tri 23703 34505 23711 34513 sw
rect 23596 34497 23711 34505
tri 23711 34497 23719 34505 sw
rect 70802 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 23596 34489 23719 34497
tri 23719 34489 23727 34497 sw
rect 23596 34482 23727 34489
rect 23462 34481 23727 34482
tri 23727 34481 23735 34489 sw
rect 23462 34478 23735 34481
tri 23462 34470 23470 34478 ne
rect 23470 34475 23735 34478
tri 23735 34475 23741 34481 sw
rect 23470 34470 23741 34475
tri 23470 34462 23478 34470 ne
rect 23478 34467 23741 34470
tri 23741 34467 23749 34475 sw
rect 23478 34462 23749 34467
tri 23478 34454 23486 34462 ne
rect 23486 34459 23749 34462
tri 23749 34459 23757 34467 sw
rect 23486 34454 23757 34459
tri 23486 34451 23489 34454 ne
rect 23489 34451 23757 34454
tri 23757 34451 23765 34459 sw
tri 23489 34443 23497 34451 ne
rect 23497 34443 23765 34451
tri 23765 34443 23773 34451 sw
rect 70802 34444 71000 34502
tri 23497 34435 23505 34443 ne
rect 23505 34435 23773 34443
tri 23773 34435 23781 34443 sw
tri 23505 34427 23513 34435 ne
rect 23513 34427 23781 34435
tri 23781 34427 23789 34435 sw
tri 23513 34419 23521 34427 ne
rect 23521 34419 23789 34427
tri 23789 34419 23797 34427 sw
tri 23521 34411 23529 34419 ne
rect 23529 34411 23797 34419
tri 23797 34411 23805 34419 sw
tri 23529 34403 23537 34411 ne
rect 23537 34403 23805 34411
tri 23805 34403 23813 34411 sw
tri 23537 34395 23545 34403 ne
rect 23545 34396 23813 34403
rect 23545 34395 23682 34396
tri 23545 34387 23553 34395 ne
rect 23553 34387 23682 34395
tri 23553 34379 23561 34387 ne
rect 23561 34379 23682 34387
tri 23561 34371 23569 34379 ne
rect 23569 34371 23682 34379
tri 23569 34363 23577 34371 ne
rect 23577 34363 23682 34371
tri 23577 34355 23585 34363 ne
rect 23585 34355 23682 34363
tri 23585 34347 23593 34355 ne
rect 23593 34350 23682 34355
rect 23728 34395 23813 34396
tri 23813 34395 23821 34403 sw
rect 70802 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 23728 34387 23821 34395
tri 23821 34387 23829 34395 sw
rect 23728 34379 23829 34387
tri 23829 34379 23837 34387 sw
rect 23728 34371 23837 34379
tri 23837 34371 23845 34379 sw
rect 23728 34363 23845 34371
tri 23845 34363 23853 34371 sw
rect 23728 34355 23853 34363
tri 23853 34355 23861 34363 sw
rect 23728 34350 23861 34355
rect 23593 34347 23861 34350
tri 23861 34347 23869 34355 sw
tri 23593 34339 23601 34347 ne
rect 23601 34339 23869 34347
tri 23869 34339 23877 34347 sw
rect 70802 34340 71000 34398
tri 23601 34333 23607 34339 ne
rect 23607 34333 23877 34339
tri 23877 34333 23883 34339 sw
tri 23607 34325 23615 34333 ne
rect 23615 34325 23883 34333
tri 23883 34325 23891 34333 sw
tri 23615 34317 23623 34325 ne
rect 23623 34317 23891 34325
tri 23891 34317 23899 34325 sw
tri 23623 34309 23631 34317 ne
rect 23631 34309 23899 34317
tri 23899 34309 23907 34317 sw
tri 23631 34301 23639 34309 ne
rect 23639 34301 23907 34309
tri 23907 34301 23915 34309 sw
tri 23639 34293 23647 34301 ne
rect 23647 34293 23915 34301
tri 23915 34293 23923 34301 sw
rect 70802 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23647 34285 23655 34293 ne
rect 23655 34285 23923 34293
tri 23923 34285 23931 34293 sw
tri 23655 34277 23663 34285 ne
rect 23663 34277 23931 34285
tri 23931 34277 23939 34285 sw
tri 23663 34269 23671 34277 ne
rect 23671 34269 23939 34277
tri 23939 34269 23947 34277 sw
tri 23671 34261 23679 34269 ne
rect 23679 34264 23947 34269
rect 23679 34261 23814 34264
tri 23679 34253 23687 34261 ne
rect 23687 34253 23814 34261
tri 23687 34245 23695 34253 ne
rect 23695 34245 23814 34253
tri 23695 34237 23703 34245 ne
rect 23703 34237 23814 34245
tri 23703 34229 23711 34237 ne
rect 23711 34229 23814 34237
tri 23711 34221 23719 34229 ne
rect 23719 34221 23814 34229
tri 23719 34213 23727 34221 ne
rect 23727 34218 23814 34221
rect 23860 34261 23947 34264
tri 23947 34261 23955 34269 sw
rect 23860 34253 23955 34261
tri 23955 34253 23963 34261 sw
rect 23860 34245 23963 34253
tri 23963 34245 23971 34253 sw
rect 23860 34237 23971 34245
tri 23971 34237 23979 34245 sw
rect 23860 34229 23979 34237
tri 23979 34229 23987 34237 sw
rect 70802 34236 71000 34294
rect 23860 34227 23987 34229
tri 23987 34227 23989 34229 sw
rect 23860 34219 23989 34227
tri 23989 34219 23997 34227 sw
rect 23860 34218 23997 34219
rect 23727 34213 23997 34218
tri 23727 34210 23730 34213 ne
rect 23730 34211 23997 34213
tri 23997 34211 24005 34219 sw
rect 23730 34210 24005 34211
tri 23730 34202 23738 34210 ne
rect 23738 34203 24005 34210
tri 24005 34203 24013 34211 sw
rect 23738 34202 24013 34203
tri 23738 34194 23746 34202 ne
rect 23746 34195 24013 34202
tri 24013 34195 24021 34203 sw
rect 23746 34194 24021 34195
tri 23746 34186 23754 34194 ne
rect 23754 34187 24021 34194
tri 24021 34187 24029 34195 sw
rect 70802 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 23754 34186 24029 34187
tri 23754 34178 23762 34186 ne
rect 23762 34179 24029 34186
tri 24029 34179 24037 34187 sw
rect 23762 34178 24037 34179
tri 23762 34170 23770 34178 ne
rect 23770 34171 24037 34178
tri 24037 34171 24045 34179 sw
rect 23770 34170 24045 34171
tri 23770 34162 23778 34170 ne
rect 23778 34163 24045 34170
tri 24045 34163 24053 34171 sw
rect 23778 34162 24053 34163
tri 23778 34154 23786 34162 ne
rect 23786 34159 24053 34162
tri 24053 34159 24057 34163 sw
rect 23786 34154 24057 34159
tri 23786 34146 23794 34154 ne
rect 23794 34151 24057 34154
tri 24057 34151 24065 34159 sw
rect 23794 34146 24065 34151
tri 23794 34138 23802 34146 ne
rect 23802 34143 24065 34146
tri 24065 34143 24073 34151 sw
rect 23802 34138 24073 34143
tri 23802 34130 23810 34138 ne
rect 23810 34135 24073 34138
tri 24073 34135 24081 34143 sw
rect 23810 34132 24081 34135
rect 23810 34130 23946 34132
tri 23810 34122 23818 34130 ne
rect 23818 34122 23946 34130
tri 23818 34114 23826 34122 ne
rect 23826 34114 23946 34122
tri 23826 34106 23834 34114 ne
rect 23834 34106 23946 34114
tri 23834 34098 23842 34106 ne
rect 23842 34098 23946 34106
tri 23842 34090 23850 34098 ne
rect 23850 34090 23946 34098
tri 23850 34082 23858 34090 ne
rect 23858 34086 23946 34090
rect 23992 34130 24081 34132
tri 24081 34130 24086 34135 sw
rect 70802 34132 71000 34190
rect 23992 34122 24086 34130
tri 24086 34122 24094 34130 sw
rect 23992 34114 24094 34122
tri 24094 34114 24102 34122 sw
rect 23992 34106 24102 34114
tri 24102 34106 24110 34114 sw
rect 23992 34098 24110 34106
tri 24110 34098 24118 34106 sw
rect 23992 34090 24118 34098
tri 24118 34090 24126 34098 sw
rect 23992 34086 24126 34090
rect 23858 34082 24126 34086
tri 24126 34082 24134 34090 sw
rect 70802 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
tri 23858 34074 23866 34082 ne
rect 23866 34074 24134 34082
tri 24134 34074 24142 34082 sw
tri 23866 34068 23872 34074 ne
rect 23872 34073 24142 34074
tri 24142 34073 24143 34074 sw
rect 23872 34068 24143 34073
tri 23872 34060 23880 34068 ne
rect 23880 34065 24143 34068
tri 24143 34065 24151 34073 sw
rect 23880 34060 24151 34065
tri 23880 34052 23888 34060 ne
rect 23888 34057 24151 34060
tri 24151 34057 24159 34065 sw
rect 23888 34052 24159 34057
tri 23888 34044 23896 34052 ne
rect 23896 34049 24159 34052
tri 24159 34049 24167 34057 sw
rect 23896 34044 24167 34049
tri 23896 34036 23904 34044 ne
rect 23904 34041 24167 34044
tri 24167 34041 24175 34049 sw
rect 23904 34036 24175 34041
tri 23904 34028 23912 34036 ne
rect 23912 34033 24175 34036
tri 24175 34033 24183 34041 sw
rect 23912 34028 24183 34033
tri 23912 34020 23920 34028 ne
rect 23920 34025 24183 34028
tri 24183 34025 24191 34033 sw
rect 70802 34028 71000 34086
rect 23920 34020 24191 34025
tri 23920 34012 23928 34020 ne
rect 23928 34017 24191 34020
tri 24191 34017 24199 34025 sw
rect 23928 34012 24199 34017
tri 23928 34004 23936 34012 ne
rect 23936 34009 24199 34012
tri 24199 34009 24207 34017 sw
rect 23936 34004 24207 34009
tri 23936 33996 23944 34004 ne
rect 23944 34001 24207 34004
tri 24207 34001 24215 34009 sw
rect 23944 34000 24215 34001
rect 23944 33996 24078 34000
tri 23944 33988 23952 33996 ne
rect 23952 33988 24078 33996
tri 23952 33980 23960 33988 ne
rect 23960 33980 24078 33988
tri 23960 33975 23965 33980 ne
rect 23965 33975 24078 33980
tri 23965 33967 23973 33975 ne
rect 23973 33967 24078 33975
tri 23973 33959 23981 33967 ne
rect 23981 33959 24078 33967
tri 23981 33951 23989 33959 ne
rect 23989 33954 24078 33959
rect 24124 33993 24215 34000
tri 24215 33993 24223 34001 sw
rect 24124 33985 24223 33993
tri 24223 33985 24231 33993 sw
rect 24124 33977 24231 33985
tri 24231 33977 24239 33985 sw
rect 70802 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33969 24239 33977
tri 24239 33969 24247 33977 sw
rect 24124 33961 24247 33969
tri 24247 33961 24255 33969 sw
rect 24124 33954 24255 33961
rect 23989 33953 24255 33954
tri 24255 33953 24263 33961 sw
rect 23989 33951 24263 33953
tri 23989 33943 23997 33951 ne
rect 23997 33945 24263 33951
tri 24263 33945 24271 33953 sw
rect 23997 33943 24271 33945
tri 23997 33935 24005 33943 ne
rect 24005 33939 24271 33943
tri 24271 33939 24277 33945 sw
rect 24005 33935 24277 33939
tri 24005 33927 24013 33935 ne
rect 24013 33931 24277 33935
tri 24277 33931 24285 33939 sw
rect 24013 33927 24285 33931
tri 24013 33919 24021 33927 ne
rect 24021 33923 24285 33927
tri 24285 33923 24293 33931 sw
rect 70802 33924 71000 33982
rect 24021 33919 24293 33923
tri 24021 33911 24029 33919 ne
rect 24029 33915 24293 33919
tri 24293 33915 24301 33923 sw
rect 24029 33911 24301 33915
tri 24029 33903 24037 33911 ne
rect 24037 33907 24301 33911
tri 24301 33907 24309 33915 sw
rect 24037 33903 24309 33907
tri 24037 33895 24045 33903 ne
rect 24045 33899 24309 33903
tri 24309 33899 24317 33907 sw
rect 24045 33895 24317 33899
tri 24045 33891 24049 33895 ne
rect 24049 33891 24317 33895
tri 24317 33891 24325 33899 sw
tri 24049 33883 24057 33891 ne
rect 24057 33883 24325 33891
tri 24325 33883 24333 33891 sw
tri 24057 33875 24065 33883 ne
rect 24065 33875 24333 33883
tri 24333 33875 24341 33883 sw
rect 70802 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
tri 24065 33867 24073 33875 ne
rect 24073 33868 24341 33875
rect 24073 33867 24210 33868
tri 24073 33859 24081 33867 ne
rect 24081 33859 24210 33867
tri 24081 33851 24089 33859 ne
rect 24089 33851 24210 33859
tri 24089 33843 24097 33851 ne
rect 24097 33843 24210 33851
tri 24097 33835 24105 33843 ne
rect 24105 33835 24210 33843
tri 24105 33827 24113 33835 ne
rect 24113 33827 24210 33835
tri 24113 33819 24121 33827 ne
rect 24121 33822 24210 33827
rect 24256 33867 24341 33868
tri 24341 33867 24349 33875 sw
rect 24256 33859 24349 33867
tri 24349 33859 24357 33867 sw
rect 24256 33851 24357 33859
tri 24357 33851 24365 33859 sw
rect 24256 33843 24365 33851
tri 24365 33843 24373 33851 sw
rect 24256 33835 24373 33843
tri 24373 33835 24381 33843 sw
rect 24256 33827 24381 33835
tri 24381 33827 24389 33835 sw
rect 24256 33822 24389 33827
rect 24121 33819 24389 33822
tri 24389 33819 24397 33827 sw
rect 70802 33820 71000 33878
tri 24121 33811 24129 33819 ne
rect 24129 33811 24397 33819
tri 24397 33811 24405 33819 sw
tri 24129 33803 24137 33811 ne
rect 24137 33803 24405 33811
tri 24405 33803 24413 33811 sw
tri 24137 33800 24140 33803 ne
rect 24140 33800 24413 33803
tri 24413 33800 24416 33803 sw
tri 24140 33792 24148 33800 ne
rect 24148 33792 24416 33800
tri 24416 33792 24424 33800 sw
tri 24148 33784 24156 33792 ne
rect 24156 33784 24424 33792
tri 24424 33784 24432 33792 sw
tri 24156 33776 24164 33784 ne
rect 24164 33776 24432 33784
tri 24432 33776 24440 33784 sw
tri 24164 33768 24172 33776 ne
rect 24172 33768 24440 33776
tri 24440 33768 24448 33776 sw
rect 70802 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24172 33760 24180 33768 ne
rect 24180 33760 24448 33768
tri 24448 33760 24456 33768 sw
tri 24180 33752 24188 33760 ne
rect 24188 33752 24456 33760
tri 24456 33752 24464 33760 sw
tri 24188 33744 24196 33752 ne
rect 24196 33744 24464 33752
tri 24464 33744 24472 33752 sw
tri 24196 33736 24204 33744 ne
rect 24204 33736 24472 33744
tri 24472 33736 24480 33744 sw
tri 24204 33728 24212 33736 ne
rect 24212 33728 24342 33736
tri 24212 33720 24220 33728 ne
rect 24220 33720 24342 33728
tri 24220 33712 24228 33720 ne
rect 24228 33712 24342 33720
tri 24228 33704 24236 33712 ne
rect 24236 33704 24342 33712
tri 24236 33696 24244 33704 ne
rect 24244 33696 24342 33704
tri 24244 33688 24252 33696 ne
rect 24252 33690 24342 33696
rect 24388 33728 24480 33736
tri 24480 33728 24488 33736 sw
rect 24388 33720 24488 33728
tri 24488 33720 24496 33728 sw
rect 24388 33712 24496 33720
tri 24496 33712 24504 33720 sw
rect 70802 33716 71000 33774
rect 24388 33704 24504 33712
tri 24504 33704 24512 33712 sw
rect 24388 33696 24512 33704
tri 24512 33696 24520 33704 sw
rect 24388 33690 24520 33696
rect 24252 33688 24520 33690
tri 24520 33688 24528 33696 sw
tri 24252 33680 24260 33688 ne
rect 24260 33682 24528 33688
tri 24528 33682 24534 33688 sw
rect 24260 33680 24534 33682
tri 24260 33674 24266 33680 ne
rect 24266 33674 24534 33680
tri 24534 33674 24542 33682 sw
tri 24266 33666 24274 33674 ne
rect 24274 33666 24542 33674
tri 24542 33666 24550 33674 sw
rect 70802 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
tri 24274 33658 24282 33666 ne
rect 24282 33658 24550 33666
tri 24550 33658 24558 33666 sw
tri 24282 33650 24290 33658 ne
rect 24290 33650 24558 33658
tri 24558 33650 24566 33658 sw
tri 24290 33642 24298 33650 ne
rect 24298 33642 24566 33650
tri 24566 33642 24574 33650 sw
tri 24298 33634 24306 33642 ne
rect 24306 33634 24574 33642
tri 24574 33634 24582 33642 sw
tri 24306 33626 24314 33634 ne
rect 24314 33626 24582 33634
tri 24582 33626 24590 33634 sw
tri 24314 33618 24322 33626 ne
rect 24322 33618 24590 33626
tri 24590 33618 24598 33626 sw
tri 24322 33610 24330 33618 ne
rect 24330 33610 24598 33618
tri 24598 33610 24606 33618 sw
rect 70802 33612 71000 33670
tri 24330 33602 24338 33610 ne
rect 24338 33604 24606 33610
rect 24338 33602 24474 33604
tri 24338 33594 24346 33602 ne
rect 24346 33594 24474 33602
tri 24346 33586 24354 33594 ne
rect 24354 33586 24474 33594
tri 24354 33578 24362 33586 ne
rect 24362 33578 24474 33586
tri 24362 33570 24370 33578 ne
rect 24370 33570 24474 33578
tri 24370 33562 24378 33570 ne
rect 24378 33562 24474 33570
tri 24378 33554 24386 33562 ne
rect 24386 33558 24474 33562
rect 24520 33602 24606 33604
tri 24606 33602 24614 33610 sw
rect 24520 33594 24614 33602
tri 24614 33594 24622 33602 sw
rect 24520 33586 24622 33594
tri 24622 33586 24630 33594 sw
rect 24520 33578 24630 33586
tri 24630 33578 24638 33586 sw
rect 24520 33570 24638 33578
tri 24638 33570 24646 33578 sw
rect 24520 33562 24646 33570
tri 24646 33562 24654 33570 sw
rect 70802 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 24520 33558 24654 33562
rect 24386 33556 24654 33558
tri 24654 33556 24660 33562 sw
rect 24386 33554 24660 33556
tri 24386 33546 24394 33554 ne
rect 24394 33548 24660 33554
tri 24660 33548 24668 33556 sw
rect 24394 33546 24668 33548
tri 24394 33538 24402 33546 ne
rect 24402 33540 24668 33546
tri 24668 33540 24676 33548 sw
rect 24402 33538 24676 33540
tri 24402 33532 24408 33538 ne
rect 24408 33532 24676 33538
tri 24676 33532 24684 33540 sw
tri 24408 33524 24416 33532 ne
rect 24416 33524 24684 33532
tri 24684 33524 24692 33532 sw
tri 24416 33516 24424 33524 ne
rect 24424 33516 24692 33524
tri 24692 33516 24700 33524 sw
tri 24424 33508 24432 33516 ne
rect 24432 33508 24700 33516
tri 24700 33508 24708 33516 sw
rect 70802 33508 71000 33566
tri 24432 33500 24440 33508 ne
rect 24440 33500 24708 33508
tri 24708 33500 24716 33508 sw
tri 24440 33492 24448 33500 ne
rect 24448 33492 24716 33500
tri 24716 33492 24724 33500 sw
tri 24448 33484 24456 33492 ne
rect 24456 33484 24724 33492
tri 24724 33484 24732 33492 sw
tri 24456 33476 24464 33484 ne
rect 24464 33476 24732 33484
tri 24732 33476 24740 33484 sw
tri 24464 33468 24472 33476 ne
rect 24472 33472 24740 33476
rect 24472 33468 24606 33472
tri 24472 33460 24480 33468 ne
rect 24480 33460 24606 33468
tri 24480 33452 24488 33460 ne
rect 24488 33452 24606 33460
tri 24488 33444 24496 33452 ne
rect 24496 33444 24606 33452
tri 24496 33436 24504 33444 ne
rect 24504 33436 24606 33444
tri 24504 33428 24512 33436 ne
rect 24512 33428 24606 33436
tri 24512 33420 24520 33428 ne
rect 24520 33426 24606 33428
rect 24652 33468 24740 33472
tri 24740 33468 24748 33476 sw
rect 24652 33460 24748 33468
tri 24748 33460 24756 33468 sw
rect 70802 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24652 33452 24756 33460
tri 24756 33452 24764 33460 sw
rect 24652 33444 24764 33452
tri 24764 33444 24772 33452 sw
rect 24652 33436 24772 33444
tri 24772 33436 24780 33444 sw
rect 24652 33428 24780 33436
tri 24780 33428 24788 33436 sw
rect 24652 33426 24788 33428
rect 24520 33420 24788 33426
tri 24788 33420 24796 33428 sw
tri 24520 33412 24528 33420 ne
rect 24528 33415 24796 33420
tri 24796 33415 24801 33420 sw
rect 24528 33412 24801 33415
tri 24528 33404 24536 33412 ne
rect 24536 33407 24801 33412
tri 24801 33407 24809 33415 sw
rect 24536 33404 24809 33407
tri 24536 33399 24541 33404 ne
rect 24541 33399 24809 33404
tri 24809 33399 24817 33407 sw
rect 70802 33404 71000 33462
tri 24541 33391 24549 33399 ne
rect 24549 33391 24817 33399
tri 24817 33391 24825 33399 sw
tri 24549 33383 24557 33391 ne
rect 24557 33383 24825 33391
tri 24825 33383 24833 33391 sw
tri 24557 33375 24565 33383 ne
rect 24565 33375 24833 33383
tri 24833 33375 24841 33383 sw
tri 24565 33367 24573 33375 ne
rect 24573 33367 24841 33375
tri 24841 33367 24849 33375 sw
tri 24573 33359 24581 33367 ne
rect 24581 33359 24849 33367
tri 24849 33359 24857 33367 sw
tri 24581 33351 24589 33359 ne
rect 24589 33351 24857 33359
tri 24857 33351 24865 33359 sw
rect 70802 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
tri 24589 33343 24597 33351 ne
rect 24597 33343 24865 33351
tri 24865 33343 24873 33351 sw
tri 24597 33335 24605 33343 ne
rect 24605 33340 24873 33343
rect 24605 33335 24738 33340
tri 24605 33327 24613 33335 ne
rect 24613 33327 24738 33335
tri 24613 33326 24614 33327 ne
rect 24614 33326 24738 33327
tri 24614 33319 24621 33326 ne
rect 24621 33319 24738 33326
tri 24621 33311 24629 33319 ne
rect 24629 33311 24738 33319
tri 24629 33303 24637 33311 ne
rect 24637 33303 24738 33311
tri 24637 33295 24645 33303 ne
rect 24645 33295 24738 33303
tri 24645 33287 24653 33295 ne
rect 24653 33294 24738 33295
rect 24784 33335 24873 33340
tri 24873 33335 24881 33343 sw
rect 24784 33327 24881 33335
tri 24881 33327 24889 33335 sw
rect 24784 33319 24889 33327
tri 24889 33319 24897 33327 sw
rect 24784 33311 24897 33319
tri 24897 33311 24905 33319 sw
rect 24784 33303 24905 33311
tri 24905 33303 24913 33311 sw
rect 24784 33295 24913 33303
tri 24913 33295 24921 33303 sw
rect 70802 33300 71000 33358
rect 24784 33294 24921 33295
rect 24653 33287 24921 33294
tri 24921 33287 24929 33295 sw
tri 24653 33279 24661 33287 ne
rect 24661 33279 24929 33287
tri 24929 33279 24937 33287 sw
tri 24661 33272 24668 33279 ne
rect 24668 33272 24937 33279
tri 24937 33272 24944 33279 sw
tri 24668 33264 24676 33272 ne
rect 24676 33264 24944 33272
tri 24944 33264 24952 33272 sw
tri 24676 33256 24684 33264 ne
rect 24684 33256 24952 33264
tri 24952 33256 24960 33264 sw
tri 24684 33248 24692 33256 ne
rect 24692 33248 24960 33256
tri 24960 33248 24968 33256 sw
rect 70802 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24692 33240 24700 33248 ne
rect 24700 33240 24968 33248
tri 24968 33240 24976 33248 sw
tri 24700 33232 24708 33240 ne
rect 24708 33232 24976 33240
tri 24976 33232 24984 33240 sw
tri 24708 33224 24716 33232 ne
rect 24716 33224 24984 33232
tri 24984 33224 24992 33232 sw
tri 24716 33216 24724 33224 ne
rect 24724 33216 24992 33224
tri 24992 33216 25000 33224 sw
tri 24724 33208 24732 33216 ne
rect 24732 33208 25000 33216
tri 25000 33208 25008 33216 sw
tri 24732 33200 24740 33208 ne
rect 24740 33200 24870 33208
tri 24740 33192 24748 33200 ne
rect 24748 33192 24870 33200
tri 24748 33184 24756 33192 ne
rect 24756 33184 24870 33192
tri 24756 33176 24764 33184 ne
rect 24764 33176 24870 33184
tri 24764 33172 24768 33176 ne
rect 24768 33172 24870 33176
tri 24768 33164 24776 33172 ne
rect 24776 33164 24870 33172
tri 24776 33156 24784 33164 ne
rect 24784 33162 24870 33164
rect 24916 33200 25008 33208
tri 25008 33200 25016 33208 sw
rect 24916 33192 25016 33200
tri 25016 33192 25024 33200 sw
rect 70802 33196 71000 33254
rect 24916 33184 25024 33192
tri 25024 33184 25032 33192 sw
rect 24916 33176 25032 33184
tri 25032 33176 25040 33184 sw
rect 24916 33172 25040 33176
tri 25040 33172 25044 33176 sw
rect 24916 33164 25044 33172
tri 25044 33164 25052 33172 sw
rect 24916 33162 25052 33164
rect 24784 33156 25052 33162
tri 25052 33156 25060 33164 sw
tri 24784 33148 24792 33156 ne
rect 24792 33148 25060 33156
tri 25060 33148 25068 33156 sw
rect 70802 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
tri 24792 33140 24800 33148 ne
rect 24800 33140 25068 33148
tri 25068 33140 25076 33148 sw
tri 24800 33132 24808 33140 ne
rect 24808 33132 25076 33140
tri 25076 33132 25084 33140 sw
tri 24808 33124 24816 33132 ne
rect 24816 33124 25084 33132
tri 25084 33124 25092 33132 sw
tri 24816 33116 24824 33124 ne
rect 24824 33116 25092 33124
tri 25092 33116 25100 33124 sw
tri 24824 33108 24832 33116 ne
rect 24832 33108 25100 33116
tri 25100 33108 25108 33116 sw
tri 24832 33100 24840 33108 ne
rect 24840 33103 25108 33108
tri 25108 33103 25113 33108 sw
rect 24840 33100 25113 33103
tri 25113 33100 25116 33103 sw
tri 24840 33092 24848 33100 ne
rect 24848 33092 25116 33100
tri 25116 33092 25124 33100 sw
rect 70802 33092 71000 33150
tri 24848 33084 24856 33092 ne
rect 24856 33084 25124 33092
tri 25124 33084 25132 33092 sw
tri 24856 33076 24864 33084 ne
rect 24864 33076 25132 33084
tri 25132 33076 25140 33084 sw
tri 24864 33068 24872 33076 ne
rect 24872 33068 25002 33076
tri 24872 33060 24880 33068 ne
rect 24880 33060 25002 33068
tri 24880 33052 24888 33060 ne
rect 24888 33052 25002 33060
tri 24888 33044 24896 33052 ne
rect 24896 33044 25002 33052
tri 24896 33036 24904 33044 ne
rect 24904 33036 25002 33044
tri 24904 33033 24907 33036 ne
rect 24907 33033 25002 33036
tri 24907 33025 24915 33033 ne
rect 24915 33030 25002 33033
rect 25048 33068 25140 33076
tri 25140 33068 25148 33076 sw
rect 25048 33060 25148 33068
tri 25148 33060 25156 33068 sw
rect 25048 33052 25156 33060
tri 25156 33052 25164 33060 sw
rect 25048 33044 25164 33052
tri 25164 33044 25172 33052 sw
rect 70802 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 25048 33036 25172 33044
tri 25172 33036 25180 33044 sw
rect 25048 33033 25180 33036
tri 25180 33033 25183 33036 sw
rect 25048 33030 25183 33033
rect 24915 33025 25183 33030
tri 25183 33025 25191 33033 sw
tri 24915 33017 24923 33025 ne
rect 24923 33017 25191 33025
tri 25191 33017 25199 33025 sw
tri 24923 33009 24931 33017 ne
rect 24931 33009 25199 33017
tri 25199 33009 25207 33017 sw
tri 24931 33001 24939 33009 ne
rect 24939 33001 25207 33009
tri 25207 33001 25215 33009 sw
tri 24939 32993 24947 33001 ne
rect 24947 32993 25215 33001
tri 25215 32993 25223 33001 sw
tri 24947 32985 24955 32993 ne
rect 24955 32985 25223 32993
tri 25223 32985 25231 32993 sw
rect 70802 32988 71000 33046
tri 24955 32977 24963 32985 ne
rect 24963 32977 25231 32985
tri 25231 32977 25239 32985 sw
tri 24963 32969 24971 32977 ne
rect 24971 32969 25239 32977
tri 25239 32969 25247 32977 sw
tri 24971 32961 24979 32969 ne
rect 24979 32961 25247 32969
tri 25247 32961 25255 32969 sw
tri 24979 32953 24987 32961 ne
rect 24987 32953 25255 32961
tri 25255 32953 25263 32961 sw
tri 24987 32945 24995 32953 ne
rect 24995 32945 25263 32953
tri 25263 32945 25271 32953 sw
tri 24995 32937 25003 32945 ne
rect 25003 32944 25271 32945
rect 25003 32937 25134 32944
tri 25003 32929 25011 32937 ne
rect 25011 32929 25134 32937
tri 25011 32921 25019 32929 ne
rect 25019 32921 25134 32929
tri 25019 32913 25027 32921 ne
rect 25027 32913 25134 32921
tri 25027 32905 25035 32913 ne
rect 25035 32905 25134 32913
tri 25035 32897 25043 32905 ne
rect 25043 32898 25134 32905
rect 25180 32937 25271 32944
tri 25271 32937 25279 32945 sw
rect 70802 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32929 25279 32937
tri 25279 32929 25287 32937 sw
rect 25180 32921 25287 32929
tri 25287 32921 25295 32929 sw
rect 25180 32913 25295 32921
tri 25295 32913 25303 32921 sw
rect 25180 32905 25303 32913
tri 25303 32905 25311 32913 sw
rect 25180 32898 25311 32905
rect 25043 32897 25311 32898
tri 25311 32897 25319 32905 sw
tri 25043 32891 25049 32897 ne
rect 25049 32891 25319 32897
tri 25319 32891 25325 32897 sw
tri 25049 32883 25057 32891 ne
rect 25057 32883 25325 32891
tri 25325 32883 25333 32891 sw
rect 70802 32884 71000 32942
tri 25057 32875 25065 32883 ne
rect 25065 32875 25333 32883
tri 25333 32875 25341 32883 sw
tri 25065 32867 25073 32875 ne
rect 25073 32867 25341 32875
tri 25341 32867 25349 32875 sw
tri 25073 32859 25081 32867 ne
rect 25081 32859 25349 32867
tri 25349 32859 25357 32867 sw
tri 25081 32851 25089 32859 ne
rect 25089 32851 25357 32859
tri 25357 32851 25365 32859 sw
tri 25089 32843 25097 32851 ne
rect 25097 32843 25365 32851
tri 25365 32843 25373 32851 sw
tri 25097 32835 25105 32843 ne
rect 25105 32835 25373 32843
tri 25373 32835 25381 32843 sw
rect 70802 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
tri 25105 32827 25113 32835 ne
rect 25113 32827 25381 32835
tri 25381 32827 25389 32835 sw
tri 25113 32824 25116 32827 ne
rect 25116 32824 25389 32827
tri 25116 32819 25121 32824 ne
rect 25121 32819 25389 32824
tri 25389 32819 25397 32827 sw
tri 25121 32811 25129 32819 ne
rect 25129 32812 25397 32819
rect 25129 32811 25266 32812
tri 25129 32803 25137 32811 ne
rect 25137 32803 25266 32811
tri 25137 32795 25145 32803 ne
rect 25145 32795 25266 32803
tri 25145 32787 25153 32795 ne
rect 25153 32787 25266 32795
tri 25153 32779 25161 32787 ne
rect 25161 32779 25266 32787
tri 25161 32771 25169 32779 ne
rect 25169 32771 25266 32779
tri 25169 32763 25177 32771 ne
rect 25177 32766 25266 32771
rect 25312 32811 25397 32812
tri 25397 32811 25405 32819 sw
rect 25312 32803 25405 32811
tri 25405 32803 25413 32811 sw
rect 25312 32795 25413 32803
tri 25413 32795 25421 32803 sw
rect 25312 32787 25421 32795
tri 25421 32787 25429 32795 sw
rect 25312 32779 25429 32787
tri 25429 32779 25437 32787 sw
rect 70802 32780 71000 32838
rect 25312 32771 25437 32779
tri 25437 32771 25445 32779 sw
rect 25312 32766 25445 32771
rect 25177 32763 25445 32766
tri 25445 32763 25453 32771 sw
tri 25177 32755 25185 32763 ne
rect 25185 32755 25453 32763
tri 25453 32755 25461 32763 sw
tri 25185 32749 25191 32755 ne
rect 25191 32749 25461 32755
tri 25461 32749 25467 32755 sw
tri 25191 32741 25199 32749 ne
rect 25199 32741 25467 32749
tri 25467 32741 25475 32749 sw
tri 25199 32733 25207 32741 ne
rect 25207 32733 25475 32741
tri 25475 32733 25483 32741 sw
rect 70802 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25207 32725 25215 32733 ne
rect 25215 32725 25483 32733
tri 25483 32725 25491 32733 sw
tri 25215 32717 25223 32725 ne
rect 25223 32717 25491 32725
tri 25491 32717 25499 32725 sw
tri 25223 32709 25231 32717 ne
rect 25231 32709 25499 32717
tri 25499 32709 25507 32717 sw
tri 25231 32701 25239 32709 ne
rect 25239 32701 25507 32709
tri 25507 32701 25515 32709 sw
tri 25239 32693 25247 32701 ne
rect 25247 32693 25515 32701
tri 25515 32693 25523 32701 sw
tri 25247 32685 25255 32693 ne
rect 25255 32685 25523 32693
tri 25523 32685 25531 32693 sw
tri 25255 32677 25263 32685 ne
rect 25263 32680 25531 32685
rect 25263 32677 25398 32680
tri 25263 32669 25271 32677 ne
rect 25271 32669 25398 32677
tri 25271 32661 25279 32669 ne
rect 25279 32661 25398 32669
tri 25279 32653 25287 32661 ne
rect 25287 32653 25398 32661
tri 25287 32645 25295 32653 ne
rect 25295 32645 25398 32653
tri 25295 32637 25303 32645 ne
rect 25303 32637 25398 32645
tri 25303 32629 25311 32637 ne
rect 25311 32634 25398 32637
rect 25444 32677 25531 32680
tri 25531 32677 25539 32685 sw
rect 25444 32669 25539 32677
tri 25539 32669 25547 32677 sw
rect 70802 32676 71000 32734
rect 25444 32661 25547 32669
tri 25547 32661 25555 32669 sw
rect 25444 32653 25555 32661
tri 25555 32653 25563 32661 sw
rect 25444 32645 25563 32653
tri 25563 32645 25571 32653 sw
rect 25444 32637 25571 32645
tri 25571 32637 25579 32645 sw
rect 25444 32634 25579 32637
rect 25311 32629 25579 32634
tri 25579 32629 25587 32637 sw
rect 70802 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25311 32626 25314 32629 ne
rect 25314 32626 25587 32629
tri 25314 32618 25322 32626 ne
rect 25322 32621 25587 32626
tri 25587 32621 25595 32629 sw
rect 25322 32618 25595 32621
tri 25322 32610 25330 32618 ne
rect 25330 32613 25595 32618
tri 25595 32613 25603 32621 sw
rect 25330 32610 25603 32613
tri 25330 32602 25338 32610 ne
rect 25338 32605 25603 32610
tri 25603 32605 25611 32613 sw
rect 25338 32602 25611 32605
tri 25338 32594 25346 32602 ne
rect 25346 32597 25611 32602
tri 25611 32597 25619 32605 sw
rect 25346 32594 25619 32597
tri 25346 32586 25354 32594 ne
rect 25354 32589 25619 32594
tri 25619 32589 25627 32597 sw
rect 25354 32586 25627 32589
tri 25354 32578 25362 32586 ne
rect 25362 32581 25627 32586
tri 25627 32581 25635 32589 sw
rect 25362 32578 25635 32581
tri 25362 32570 25370 32578 ne
rect 25370 32573 25635 32578
tri 25635 32573 25643 32581 sw
rect 25370 32570 25643 32573
tri 25370 32562 25378 32570 ne
rect 25378 32565 25643 32570
tri 25643 32565 25651 32573 sw
rect 70802 32572 71000 32630
rect 25378 32562 25651 32565
tri 25378 32554 25386 32562 ne
rect 25386 32557 25651 32562
tri 25651 32557 25659 32565 sw
rect 25386 32554 25659 32557
tri 25386 32546 25394 32554 ne
rect 25394 32549 25659 32554
tri 25659 32549 25667 32557 sw
rect 25394 32548 25667 32549
rect 25394 32546 25530 32548
tri 25394 32538 25402 32546 ne
rect 25402 32538 25530 32546
tri 25402 32530 25410 32538 ne
rect 25410 32530 25530 32538
tri 25410 32522 25418 32530 ne
rect 25418 32522 25530 32530
tri 25418 32514 25426 32522 ne
rect 25426 32514 25530 32522
tri 25426 32506 25434 32514 ne
rect 25434 32506 25530 32514
tri 25434 32498 25442 32506 ne
rect 25442 32502 25530 32506
rect 25576 32541 25667 32548
tri 25667 32541 25675 32549 sw
rect 25576 32533 25675 32541
tri 25675 32533 25683 32541 sw
rect 25576 32525 25683 32533
tri 25683 32525 25691 32533 sw
rect 70802 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 25576 32517 25691 32525
tri 25691 32517 25699 32525 sw
rect 25576 32509 25699 32517
tri 25699 32509 25707 32517 sw
rect 25576 32502 25707 32509
rect 25442 32501 25707 32502
tri 25707 32501 25715 32509 sw
rect 25442 32498 25715 32501
tri 25442 32490 25450 32498 ne
rect 25450 32493 25715 32498
tri 25715 32493 25723 32501 sw
rect 25450 32490 25723 32493
tri 25450 32482 25458 32490 ne
rect 25458 32485 25723 32490
tri 25723 32485 25731 32493 sw
rect 25458 32482 25731 32485
tri 25458 32481 25459 32482 ne
rect 25459 32481 25731 32482
tri 25731 32481 25735 32485 sw
tri 25459 32473 25467 32481 ne
rect 25467 32473 25735 32481
tri 25735 32473 25743 32481 sw
tri 25467 32465 25475 32473 ne
rect 25475 32465 25743 32473
tri 25743 32465 25751 32473 sw
rect 70802 32468 71000 32526
tri 25475 32457 25483 32465 ne
rect 25483 32457 25751 32465
tri 25751 32457 25759 32465 sw
tri 25483 32449 25491 32457 ne
rect 25491 32449 25759 32457
tri 25759 32449 25767 32457 sw
tri 25491 32441 25499 32449 ne
rect 25499 32441 25767 32449
tri 25767 32441 25775 32449 sw
tri 25499 32433 25507 32441 ne
rect 25507 32433 25775 32441
tri 25775 32433 25783 32441 sw
tri 25507 32425 25515 32433 ne
rect 25515 32425 25783 32433
tri 25783 32425 25791 32433 sw
tri 25515 32417 25523 32425 ne
rect 25523 32417 25791 32425
tri 25791 32417 25799 32425 sw
rect 70802 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
tri 25523 32409 25531 32417 ne
rect 25531 32416 25799 32417
rect 25531 32409 25662 32416
tri 25531 32401 25539 32409 ne
rect 25539 32401 25662 32409
tri 25539 32393 25547 32401 ne
rect 25547 32393 25662 32401
tri 25547 32385 25555 32393 ne
rect 25555 32385 25662 32393
tri 25555 32377 25563 32385 ne
rect 25563 32377 25662 32385
tri 25563 32369 25571 32377 ne
rect 25571 32370 25662 32377
rect 25708 32409 25799 32416
tri 25799 32409 25807 32417 sw
rect 25708 32401 25807 32409
tri 25807 32401 25815 32409 sw
rect 25708 32393 25815 32401
tri 25815 32393 25823 32401 sw
rect 25708 32385 25823 32393
tri 25823 32385 25831 32393 sw
rect 25708 32377 25831 32385
tri 25831 32377 25839 32385 sw
rect 25708 32370 25839 32377
rect 25571 32369 25839 32370
tri 25839 32369 25847 32377 sw
tri 25571 32361 25579 32369 ne
rect 25579 32361 25847 32369
tri 25847 32361 25855 32369 sw
rect 70802 32364 71000 32422
tri 25579 32353 25587 32361 ne
rect 25587 32353 25855 32361
tri 25855 32353 25863 32361 sw
tri 25587 32351 25589 32353 ne
rect 25589 32351 25863 32353
tri 25863 32351 25865 32353 sw
tri 25589 32343 25597 32351 ne
rect 25597 32343 25865 32351
tri 25865 32343 25873 32351 sw
tri 25597 32335 25605 32343 ne
rect 25605 32335 25873 32343
tri 25873 32335 25881 32343 sw
tri 25605 32327 25613 32335 ne
rect 25613 32327 25881 32335
tri 25881 32327 25889 32335 sw
tri 25613 32319 25621 32327 ne
rect 25621 32319 25889 32327
tri 25889 32319 25897 32327 sw
tri 25621 32311 25629 32319 ne
rect 25629 32311 25897 32319
tri 25897 32311 25905 32319 sw
rect 70802 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
tri 25629 32303 25637 32311 ne
rect 25637 32303 25905 32311
tri 25905 32303 25913 32311 sw
tri 25637 32295 25645 32303 ne
rect 25645 32295 25913 32303
tri 25913 32295 25921 32303 sw
tri 25645 32287 25653 32295 ne
rect 25653 32287 25921 32295
tri 25921 32287 25929 32295 sw
tri 25653 32279 25661 32287 ne
rect 25661 32284 25929 32287
rect 25661 32279 25794 32284
tri 25661 32271 25669 32279 ne
rect 25669 32271 25794 32279
tri 25669 32263 25677 32271 ne
rect 25677 32263 25794 32271
tri 25677 32255 25685 32263 ne
rect 25685 32255 25794 32263
tri 25685 32247 25693 32255 ne
rect 25693 32247 25794 32255
tri 25693 32239 25701 32247 ne
rect 25701 32239 25794 32247
tri 25701 32231 25709 32239 ne
rect 25709 32238 25794 32239
rect 25840 32279 25929 32284
tri 25929 32279 25937 32287 sw
rect 25840 32271 25937 32279
tri 25937 32271 25945 32279 sw
rect 25840 32263 25945 32271
tri 25945 32263 25953 32271 sw
rect 25840 32255 25953 32263
tri 25953 32255 25961 32263 sw
rect 70802 32260 71000 32318
rect 25840 32247 25961 32255
tri 25961 32247 25969 32255 sw
rect 25840 32239 25969 32247
tri 25969 32239 25977 32247 sw
rect 25840 32238 25977 32239
rect 25709 32231 25977 32238
tri 25977 32231 25985 32239 sw
tri 25709 32223 25717 32231 ne
rect 25717 32226 25985 32231
tri 25985 32226 25990 32231 sw
rect 25717 32223 25990 32226
tri 25717 32215 25725 32223 ne
rect 25725 32218 25990 32223
tri 25990 32218 25998 32226 sw
rect 25725 32215 25998 32218
tri 25725 32210 25730 32215 ne
rect 25730 32210 25998 32215
tri 25998 32210 26006 32218 sw
rect 70802 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25730 32202 25738 32210 ne
rect 25738 32202 26006 32210
tri 26006 32202 26014 32210 sw
tri 25738 32194 25746 32202 ne
rect 25746 32194 26014 32202
tri 26014 32194 26022 32202 sw
tri 25746 32186 25754 32194 ne
rect 25754 32186 26022 32194
tri 26022 32186 26030 32194 sw
tri 25754 32178 25762 32186 ne
rect 25762 32178 26030 32186
tri 26030 32178 26038 32186 sw
tri 25762 32170 25770 32178 ne
rect 25770 32170 26038 32178
tri 26038 32170 26046 32178 sw
tri 25770 32162 25778 32170 ne
rect 25778 32162 26046 32170
tri 26046 32162 26054 32170 sw
tri 25778 32154 25786 32162 ne
rect 25786 32154 26054 32162
tri 26054 32154 26062 32162 sw
rect 70802 32156 71000 32214
tri 25786 32146 25794 32154 ne
rect 25794 32152 26062 32154
rect 25794 32146 25926 32152
tri 25794 32138 25802 32146 ne
rect 25802 32138 25926 32146
tri 25802 32130 25810 32138 ne
rect 25810 32130 25926 32138
tri 25810 32122 25818 32130 ne
rect 25818 32122 25926 32130
tri 25818 32114 25826 32122 ne
rect 25826 32114 25926 32122
tri 25826 32106 25834 32114 ne
rect 25834 32106 25926 32114
rect 25972 32146 26062 32152
tri 26062 32146 26070 32154 sw
rect 25972 32138 26070 32146
tri 26070 32138 26078 32146 sw
rect 25972 32130 26078 32138
tri 26078 32130 26086 32138 sw
rect 25972 32122 26086 32130
tri 26086 32122 26094 32130 sw
rect 25972 32116 26094 32122
tri 26094 32116 26100 32122 sw
rect 25972 32108 26100 32116
tri 26100 32108 26108 32116 sw
rect 70802 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 25972 32106 26108 32108
tri 25834 32098 25842 32106 ne
rect 25842 32100 26108 32106
tri 26108 32100 26116 32108 sw
rect 25842 32098 26116 32100
tri 25842 32090 25850 32098 ne
rect 25850 32092 26116 32098
tri 26116 32092 26124 32100 sw
rect 25850 32090 26124 32092
tri 25850 32082 25858 32090 ne
rect 25858 32084 26124 32090
tri 26124 32084 26132 32092 sw
rect 25858 32082 26132 32084
tri 25858 32074 25866 32082 ne
rect 25866 32076 26132 32082
tri 26132 32076 26140 32084 sw
rect 25866 32074 26140 32076
tri 25866 32066 25874 32074 ne
rect 25874 32068 26140 32074
tri 26140 32068 26148 32076 sw
rect 25874 32066 26148 32068
tri 25874 32058 25882 32066 ne
rect 25882 32060 26148 32066
tri 26148 32060 26156 32068 sw
rect 25882 32058 26156 32060
tri 25882 32050 25890 32058 ne
rect 25890 32052 26156 32058
tri 26156 32052 26164 32060 sw
rect 70802 32052 71000 32110
rect 25890 32050 26164 32052
tri 25890 32042 25898 32050 ne
rect 25898 32044 26164 32050
tri 26164 32044 26172 32052 sw
rect 25898 32042 26172 32044
tri 25898 32034 25906 32042 ne
rect 25906 32036 26172 32042
tri 26172 32036 26180 32044 sw
rect 25906 32034 26180 32036
tri 25906 32026 25914 32034 ne
rect 25914 32028 26180 32034
tri 26180 32028 26188 32036 sw
rect 25914 32026 26188 32028
tri 25914 32018 25922 32026 ne
rect 25922 32020 26188 32026
tri 26188 32020 26196 32028 sw
rect 25922 32018 26058 32020
tri 25922 32010 25930 32018 ne
rect 25930 32010 26058 32018
tri 25930 32003 25937 32010 ne
rect 25937 32003 26058 32010
tri 25937 31995 25945 32003 ne
rect 25945 31995 26058 32003
tri 25945 31987 25953 31995 ne
rect 25953 31987 26058 31995
tri 25953 31979 25961 31987 ne
rect 25961 31979 26058 31987
tri 25961 31971 25969 31979 ne
rect 25969 31974 26058 31979
rect 26104 32019 26196 32020
tri 26196 32019 26197 32020 sw
rect 26104 32011 26197 32019
tri 26197 32011 26205 32019 sw
rect 26104 32003 26205 32011
tri 26205 32003 26213 32011 sw
rect 70802 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 26104 31995 26213 32003
tri 26213 31995 26221 32003 sw
rect 26104 31987 26221 31995
tri 26221 31987 26229 31995 sw
rect 26104 31979 26229 31987
tri 26229 31979 26237 31987 sw
rect 26104 31974 26237 31979
rect 25969 31971 26237 31974
tri 26237 31971 26245 31979 sw
tri 25969 31963 25977 31971 ne
rect 25977 31963 26245 31971
tri 26245 31963 26253 31971 sw
tri 25977 31955 25985 31963 ne
rect 25985 31955 26253 31963
tri 26253 31955 26261 31963 sw
tri 25985 31947 25993 31955 ne
rect 25993 31947 26261 31955
tri 26261 31947 26269 31955 sw
rect 70802 31948 71000 32006
tri 25993 31939 26001 31947 ne
rect 26001 31942 26269 31947
tri 26269 31942 26274 31947 sw
rect 26001 31939 26274 31942
tri 26001 31931 26009 31939 ne
rect 26009 31934 26274 31939
tri 26274 31934 26282 31942 sw
rect 26009 31931 26282 31934
tri 26009 31930 26010 31931 ne
rect 26010 31930 26282 31931
tri 26010 31922 26018 31930 ne
rect 26018 31926 26282 31930
tri 26282 31926 26290 31934 sw
rect 26018 31922 26290 31926
tri 26018 31914 26026 31922 ne
rect 26026 31918 26290 31922
tri 26290 31918 26298 31926 sw
rect 26026 31914 26298 31918
tri 26026 31906 26034 31914 ne
rect 26034 31910 26298 31914
tri 26298 31910 26306 31918 sw
rect 26034 31906 26306 31910
tri 26034 31898 26042 31906 ne
rect 26042 31902 26306 31906
tri 26306 31902 26314 31910 sw
rect 70802 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26042 31898 26314 31902
tri 26042 31890 26050 31898 ne
rect 26050 31894 26314 31898
tri 26314 31894 26322 31902 sw
rect 26050 31890 26322 31894
tri 26050 31882 26058 31890 ne
rect 26058 31888 26322 31890
rect 26058 31882 26190 31888
tri 26058 31874 26066 31882 ne
rect 26066 31874 26190 31882
tri 26066 31866 26074 31874 ne
rect 26074 31866 26190 31874
tri 26074 31858 26082 31866 ne
rect 26082 31858 26190 31866
tri 26082 31850 26090 31858 ne
rect 26090 31850 26190 31858
tri 26090 31842 26098 31850 ne
rect 26098 31842 26190 31850
rect 26236 31886 26322 31888
tri 26322 31886 26330 31894 sw
rect 26236 31878 26330 31886
tri 26330 31878 26338 31886 sw
rect 26236 31870 26338 31878
tri 26338 31870 26346 31878 sw
rect 26236 31862 26346 31870
tri 26346 31862 26354 31870 sw
rect 26236 31854 26354 31862
tri 26354 31854 26362 31862 sw
rect 26236 31846 26362 31854
tri 26362 31846 26370 31854 sw
rect 26236 31842 26370 31846
tri 26098 31834 26106 31842 ne
rect 26106 31840 26370 31842
tri 26370 31840 26376 31846 sw
rect 70802 31844 71000 31902
rect 26106 31834 26376 31840
tri 26106 31826 26114 31834 ne
rect 26114 31832 26376 31834
tri 26376 31832 26384 31840 sw
rect 26114 31826 26384 31832
tri 26114 31823 26117 31826 ne
rect 26117 31824 26384 31826
tri 26384 31824 26392 31832 sw
rect 26117 31823 26392 31824
tri 26117 31815 26125 31823 ne
rect 26125 31816 26392 31823
tri 26392 31816 26400 31824 sw
rect 26125 31815 26400 31816
tri 26125 31807 26133 31815 ne
rect 26133 31808 26400 31815
tri 26400 31808 26408 31816 sw
rect 26133 31807 26408 31808
tri 26133 31799 26141 31807 ne
rect 26141 31800 26408 31807
tri 26408 31800 26416 31808 sw
rect 26141 31799 26416 31800
tri 26141 31791 26149 31799 ne
rect 26149 31792 26416 31799
tri 26416 31792 26424 31800 sw
rect 70802 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26149 31791 26424 31792
tri 26149 31783 26157 31791 ne
rect 26157 31784 26424 31791
tri 26424 31784 26432 31792 sw
rect 26157 31783 26432 31784
tri 26157 31775 26165 31783 ne
rect 26165 31776 26432 31783
tri 26432 31776 26440 31784 sw
rect 26165 31775 26440 31776
tri 26165 31767 26173 31775 ne
rect 26173 31768 26440 31775
tri 26440 31768 26448 31776 sw
rect 26173 31767 26448 31768
tri 26448 31767 26449 31768 sw
tri 26173 31759 26181 31767 ne
rect 26181 31759 26449 31767
tri 26449 31759 26457 31767 sw
tri 26181 31751 26189 31759 ne
rect 26189 31756 26457 31759
rect 26189 31751 26322 31756
tri 26189 31743 26197 31751 ne
rect 26197 31743 26322 31751
tri 26197 31735 26205 31743 ne
rect 26205 31735 26322 31743
tri 26205 31727 26213 31735 ne
rect 26213 31727 26322 31735
tri 26213 31719 26221 31727 ne
rect 26221 31719 26322 31727
tri 26221 31711 26229 31719 ne
rect 26229 31711 26322 31719
tri 26229 31703 26237 31711 ne
rect 26237 31710 26322 31711
rect 26368 31751 26457 31756
tri 26457 31751 26465 31759 sw
rect 26368 31743 26465 31751
tri 26465 31743 26473 31751 sw
rect 26368 31735 26473 31743
tri 26473 31735 26481 31743 sw
rect 70802 31740 71000 31798
rect 26368 31727 26481 31735
tri 26481 31727 26489 31735 sw
rect 26368 31719 26489 31727
tri 26489 31719 26497 31727 sw
rect 26368 31711 26497 31719
tri 26497 31711 26505 31719 sw
rect 26368 31710 26505 31711
rect 26237 31703 26505 31710
tri 26505 31703 26513 31711 sw
tri 26237 31695 26245 31703 ne
rect 26245 31695 26513 31703
tri 26513 31695 26521 31703 sw
tri 26245 31687 26253 31695 ne
rect 26253 31690 26521 31695
tri 26521 31690 26526 31695 sw
rect 70802 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
rect 26253 31687 26526 31690
tri 26253 31682 26258 31687 ne
rect 26258 31682 26526 31687
tri 26526 31682 26534 31690 sw
tri 26258 31674 26266 31682 ne
rect 26266 31674 26534 31682
tri 26534 31674 26542 31682 sw
tri 26266 31666 26274 31674 ne
rect 26274 31666 26542 31674
tri 26542 31666 26550 31674 sw
tri 26274 31658 26282 31666 ne
rect 26282 31658 26550 31666
tri 26550 31658 26558 31666 sw
tri 26282 31650 26290 31658 ne
rect 26290 31650 26558 31658
tri 26558 31650 26566 31658 sw
tri 26290 31642 26298 31650 ne
rect 26298 31642 26566 31650
tri 26566 31642 26574 31650 sw
tri 26298 31634 26306 31642 ne
rect 26306 31634 26574 31642
tri 26574 31634 26582 31642 sw
rect 70802 31636 71000 31694
tri 26306 31626 26314 31634 ne
rect 26314 31626 26582 31634
tri 26582 31626 26590 31634 sw
tri 26314 31618 26322 31626 ne
rect 26322 31624 26590 31626
rect 26322 31618 26454 31624
tri 26322 31610 26330 31618 ne
rect 26330 31610 26454 31618
tri 26330 31602 26338 31610 ne
rect 26338 31602 26454 31610
tri 26338 31594 26346 31602 ne
rect 26346 31594 26454 31602
tri 26346 31586 26354 31594 ne
rect 26354 31586 26454 31594
tri 26354 31578 26362 31586 ne
rect 26362 31578 26454 31586
rect 26500 31618 26590 31624
tri 26590 31618 26598 31626 sw
rect 26500 31610 26598 31618
tri 26598 31610 26606 31618 sw
rect 26500 31602 26606 31610
tri 26606 31602 26614 31610 sw
rect 26500 31594 26614 31602
tri 26614 31594 26622 31602 sw
rect 26500 31586 26622 31594
tri 26622 31586 26630 31594 sw
rect 70802 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 26500 31578 26630 31586
tri 26630 31578 26638 31586 sw
tri 26362 31570 26370 31578 ne
rect 26370 31570 26638 31578
tri 26638 31570 26646 31578 sw
tri 26370 31562 26378 31570 ne
rect 26378 31563 26646 31570
tri 26646 31563 26653 31570 sw
rect 26378 31562 26653 31563
tri 26378 31555 26385 31562 ne
rect 26385 31555 26653 31562
tri 26653 31555 26661 31563 sw
tri 26385 31547 26393 31555 ne
rect 26393 31547 26661 31555
tri 26661 31547 26669 31555 sw
tri 26393 31539 26401 31547 ne
rect 26401 31539 26669 31547
tri 26669 31539 26677 31547 sw
tri 26401 31531 26409 31539 ne
rect 26409 31531 26677 31539
tri 26677 31531 26685 31539 sw
rect 70802 31532 71000 31590
tri 26409 31523 26417 31531 ne
rect 26417 31523 26685 31531
tri 26685 31523 26693 31531 sw
tri 26417 31515 26425 31523 ne
rect 26425 31515 26693 31523
tri 26693 31515 26701 31523 sw
tri 26425 31507 26433 31515 ne
rect 26433 31507 26701 31515
tri 26701 31507 26709 31515 sw
tri 26433 31499 26441 31507 ne
rect 26441 31499 26709 31507
tri 26709 31499 26717 31507 sw
tri 26441 31491 26449 31499 ne
rect 26449 31492 26717 31499
rect 26449 31491 26586 31492
tri 26449 31483 26457 31491 ne
rect 26457 31483 26586 31491
tri 26457 31475 26465 31483 ne
rect 26465 31475 26586 31483
tri 26465 31467 26473 31475 ne
rect 26473 31467 26586 31475
tri 26473 31459 26481 31467 ne
rect 26481 31459 26586 31467
tri 26481 31451 26489 31459 ne
rect 26489 31451 26586 31459
tri 26489 31443 26497 31451 ne
rect 26497 31446 26586 31451
rect 26632 31491 26717 31492
tri 26717 31491 26725 31499 sw
rect 26632 31483 26725 31491
tri 26725 31483 26733 31491 sw
rect 70802 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31475 26733 31483
tri 26733 31475 26741 31483 sw
rect 26632 31467 26741 31475
tri 26741 31467 26749 31475 sw
rect 26632 31459 26749 31467
tri 26749 31459 26757 31467 sw
rect 26632 31451 26757 31459
tri 26757 31451 26765 31459 sw
rect 26632 31446 26765 31451
rect 26497 31443 26765 31446
tri 26765 31443 26773 31451 sw
tri 26497 31435 26505 31443 ne
rect 26505 31435 26773 31443
tri 26773 31435 26781 31443 sw
tri 26505 31427 26513 31435 ne
rect 26513 31427 26781 31435
tri 26781 31427 26789 31435 sw
rect 70802 31428 71000 31486
tri 26513 31419 26521 31427 ne
rect 26521 31419 26789 31427
tri 26789 31419 26797 31427 sw
tri 26521 31411 26529 31419 ne
rect 26529 31411 26797 31419
tri 26797 31411 26805 31419 sw
tri 26529 31403 26537 31411 ne
rect 26537 31403 26805 31411
tri 26805 31403 26813 31411 sw
tri 26537 31395 26545 31403 ne
rect 26545 31395 26813 31403
tri 26813 31395 26821 31403 sw
tri 26545 31387 26553 31395 ne
rect 26553 31387 26821 31395
tri 26821 31387 26829 31395 sw
tri 26553 31379 26561 31387 ne
rect 26561 31379 26829 31387
tri 26829 31379 26837 31387 sw
rect 70802 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
tri 26561 31371 26569 31379 ne
rect 26569 31371 26837 31379
tri 26837 31371 26845 31379 sw
tri 26569 31363 26577 31371 ne
rect 26577 31364 26845 31371
tri 26845 31364 26852 31371 sw
rect 26577 31363 26852 31364
tri 26577 31355 26585 31363 ne
rect 26585 31360 26852 31363
rect 26585 31355 26718 31360
tri 26585 31351 26589 31355 ne
rect 26589 31351 26718 31355
tri 26589 31343 26597 31351 ne
rect 26597 31343 26718 31351
tri 26597 31335 26605 31343 ne
rect 26605 31335 26718 31343
tri 26605 31327 26613 31335 ne
rect 26613 31327 26718 31335
tri 26613 31319 26621 31327 ne
rect 26621 31319 26718 31327
tri 26621 31311 26629 31319 ne
rect 26629 31314 26718 31319
rect 26764 31356 26852 31360
tri 26852 31356 26860 31364 sw
rect 26764 31348 26860 31356
tri 26860 31348 26868 31356 sw
rect 26764 31340 26868 31348
tri 26868 31340 26876 31348 sw
rect 26764 31332 26876 31340
tri 26876 31332 26884 31340 sw
rect 26764 31324 26884 31332
tri 26884 31324 26892 31332 sw
rect 70802 31324 71000 31382
rect 26764 31316 26892 31324
tri 26892 31316 26900 31324 sw
rect 26764 31314 26900 31316
rect 26629 31311 26900 31314
tri 26629 31303 26637 31311 ne
rect 26637 31308 26900 31311
tri 26900 31308 26908 31316 sw
rect 26637 31303 26908 31308
tri 26637 31295 26645 31303 ne
rect 26645 31300 26908 31303
tri 26908 31300 26916 31308 sw
rect 26645 31295 26916 31300
tri 26645 31287 26653 31295 ne
rect 26653 31292 26916 31295
tri 26916 31292 26924 31300 sw
rect 26653 31287 26924 31292
tri 26653 31279 26661 31287 ne
rect 26661 31284 26924 31287
tri 26924 31284 26932 31292 sw
rect 26661 31279 26932 31284
tri 26661 31271 26669 31279 ne
rect 26669 31276 26932 31279
tri 26932 31276 26940 31284 sw
rect 70802 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
rect 26669 31271 26940 31276
tri 26669 31263 26677 31271 ne
rect 26677 31268 26940 31271
tri 26940 31268 26948 31276 sw
rect 26677 31263 26948 31268
tri 26677 31255 26685 31263 ne
rect 26685 31260 26948 31263
tri 26948 31260 26956 31268 sw
rect 26685 31255 26956 31260
tri 26956 31255 26961 31260 sw
tri 26685 31247 26693 31255 ne
rect 26693 31247 26961 31255
tri 26961 31247 26969 31255 sw
tri 26693 31243 26697 31247 ne
rect 26697 31243 26969 31247
tri 26697 31239 26701 31243 ne
rect 26701 31239 26969 31243
tri 26969 31239 26977 31247 sw
tri 26701 31231 26709 31239 ne
rect 26709 31231 26977 31239
tri 26977 31231 26985 31239 sw
tri 26709 31223 26717 31231 ne
rect 26717 31228 26985 31231
rect 26717 31223 26850 31228
tri 26717 31215 26725 31223 ne
rect 26725 31215 26850 31223
tri 26725 31207 26733 31215 ne
rect 26733 31207 26850 31215
tri 26733 31199 26741 31207 ne
rect 26741 31199 26850 31207
tri 26741 31191 26749 31199 ne
rect 26749 31191 26850 31199
tri 26749 31183 26757 31191 ne
rect 26757 31183 26850 31191
tri 26757 31175 26765 31183 ne
rect 26765 31182 26850 31183
rect 26896 31223 26985 31228
tri 26985 31223 26993 31231 sw
rect 26896 31215 26993 31223
tri 26993 31215 27001 31223 sw
rect 70802 31220 71000 31278
rect 26896 31207 27001 31215
tri 27001 31207 27009 31215 sw
rect 26896 31199 27009 31207
tri 27009 31199 27017 31207 sw
rect 26896 31191 27017 31199
tri 27017 31191 27025 31199 sw
rect 26896 31183 27025 31191
tri 27025 31183 27033 31191 sw
rect 26896 31182 27033 31183
rect 26765 31175 27033 31182
tri 27033 31175 27041 31183 sw
tri 26765 31167 26773 31175 ne
rect 26773 31167 27041 31175
tri 27041 31167 27049 31175 sw
rect 70802 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
tri 26773 31159 26781 31167 ne
rect 26781 31159 27049 31167
tri 27049 31159 27057 31167 sw
tri 26781 31151 26789 31159 ne
rect 26789 31151 27057 31159
tri 27057 31151 27065 31159 sw
tri 26789 31143 26797 31151 ne
rect 26797 31143 27065 31151
tri 27065 31143 27073 31151 sw
tri 26797 31135 26805 31143 ne
rect 26805 31135 27073 31143
tri 27073 31135 27081 31143 sw
tri 26805 31127 26813 31135 ne
rect 26813 31127 27081 31135
tri 27081 31127 27089 31135 sw
tri 26813 31119 26821 31127 ne
rect 26821 31119 27089 31127
tri 27089 31119 27097 31127 sw
tri 26821 31111 26829 31119 ne
rect 26829 31111 27097 31119
tri 27097 31111 27105 31119 sw
rect 70802 31116 71000 31174
tri 26829 31103 26837 31111 ne
rect 26837 31103 27105 31111
tri 27105 31103 27113 31111 sw
tri 26837 31095 26845 31103 ne
rect 26845 31096 27113 31103
rect 26845 31095 26982 31096
tri 26845 31087 26853 31095 ne
rect 26853 31087 26982 31095
tri 26853 31079 26861 31087 ne
rect 26861 31079 26982 31087
tri 26861 31071 26869 31079 ne
rect 26869 31071 26982 31079
tri 26869 31063 26877 31071 ne
rect 26877 31063 26982 31071
tri 26877 31055 26885 31063 ne
rect 26885 31055 26982 31063
tri 26885 31047 26893 31055 ne
rect 26893 31050 26982 31055
rect 27028 31095 27113 31096
tri 27113 31095 27121 31103 sw
rect 27028 31087 27121 31095
tri 27121 31087 27129 31095 sw
rect 27028 31079 27129 31087
tri 27129 31079 27137 31087 sw
rect 27028 31071 27137 31079
tri 27137 31071 27145 31079 sw
rect 27028 31063 27145 31071
tri 27145 31063 27153 31071 sw
rect 70802 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 27028 31055 27153 31063
tri 27153 31055 27161 31063 sw
rect 27028 31050 27161 31055
rect 26893 31047 27161 31050
tri 27161 31047 27169 31055 sw
tri 26893 31039 26901 31047 ne
rect 26901 31039 27169 31047
tri 27169 31039 27177 31047 sw
tri 26901 31031 26909 31039 ne
rect 26909 31031 27177 31039
tri 27177 31031 27185 31039 sw
tri 26909 31023 26917 31031 ne
rect 26917 31023 27185 31031
tri 27185 31023 27193 31031 sw
tri 26917 31015 26925 31023 ne
rect 26925 31015 27193 31023
tri 27193 31015 27201 31023 sw
tri 26925 31007 26933 31015 ne
rect 26933 31007 27201 31015
tri 27201 31007 27209 31015 sw
rect 70802 31012 71000 31070
tri 26933 30999 26941 31007 ne
rect 26941 30999 27209 31007
tri 27209 30999 27217 31007 sw
tri 26941 30991 26949 30999 ne
rect 26949 30991 27217 30999
tri 27217 30991 27225 30999 sw
tri 26949 30983 26957 30991 ne
rect 26957 30983 27225 30991
tri 27225 30983 27233 30991 sw
tri 26957 30975 26965 30983 ne
rect 26965 30975 27233 30983
tri 27233 30975 27241 30983 sw
tri 26965 30971 26969 30975 ne
rect 26969 30971 27241 30975
tri 27241 30971 27245 30975 sw
tri 26969 30963 26977 30971 ne
rect 26977 30964 27245 30971
rect 26977 30963 27114 30964
tri 26977 30955 26985 30963 ne
rect 26985 30955 27114 30963
tri 26985 30947 26993 30955 ne
rect 26993 30947 27114 30955
tri 26993 30939 27001 30947 ne
rect 27001 30939 27114 30947
tri 27001 30931 27009 30939 ne
rect 27009 30931 27114 30939
tri 27009 30923 27017 30931 ne
rect 27017 30923 27114 30931
tri 27017 30915 27025 30923 ne
rect 27025 30918 27114 30923
rect 27160 30963 27245 30964
tri 27245 30963 27253 30971 sw
rect 70802 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 27160 30955 27253 30963
tri 27253 30955 27261 30963 sw
rect 27160 30947 27261 30955
tri 27261 30947 27269 30955 sw
rect 27160 30939 27269 30947
tri 27269 30939 27277 30947 sw
rect 27160 30931 27277 30939
tri 27277 30931 27285 30939 sw
rect 27160 30923 27285 30931
tri 27285 30923 27293 30931 sw
rect 27160 30918 27293 30923
rect 27025 30915 27293 30918
tri 27293 30915 27301 30923 sw
tri 27025 30907 27033 30915 ne
rect 27033 30907 27301 30915
tri 27301 30907 27309 30915 sw
rect 70802 30908 71000 30966
tri 27033 30899 27041 30907 ne
rect 27041 30899 27309 30907
tri 27309 30899 27317 30907 sw
tri 27041 30891 27049 30899 ne
rect 27049 30891 27317 30899
tri 27317 30891 27325 30899 sw
tri 27049 30883 27057 30891 ne
rect 27057 30883 27325 30891
tri 27325 30883 27333 30891 sw
tri 27057 30882 27058 30883 ne
rect 27058 30882 27333 30883
tri 27058 30874 27066 30882 ne
rect 27066 30875 27333 30882
tri 27333 30875 27341 30883 sw
rect 27066 30874 27341 30875
tri 27066 30866 27074 30874 ne
rect 27074 30867 27341 30874
tri 27341 30867 27349 30875 sw
rect 27074 30866 27349 30867
tri 27074 30858 27082 30866 ne
rect 27082 30859 27349 30866
tri 27349 30859 27357 30867 sw
rect 70802 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
rect 27082 30858 27357 30859
tri 27082 30850 27090 30858 ne
rect 27090 30851 27357 30858
tri 27357 30851 27365 30859 sw
rect 27090 30850 27365 30851
tri 27090 30842 27098 30850 ne
rect 27098 30843 27365 30850
tri 27365 30843 27373 30851 sw
rect 27098 30842 27373 30843
tri 27098 30834 27106 30842 ne
rect 27106 30835 27373 30842
tri 27373 30835 27381 30843 sw
rect 27106 30834 27381 30835
tri 27106 30826 27114 30834 ne
rect 27114 30832 27381 30834
rect 27114 30826 27246 30832
tri 27114 30818 27122 30826 ne
rect 27122 30818 27246 30826
tri 27122 30810 27130 30818 ne
rect 27130 30810 27246 30818
tri 27130 30802 27138 30810 ne
rect 27138 30802 27246 30810
tri 27138 30794 27146 30802 ne
rect 27146 30794 27246 30802
tri 27146 30786 27154 30794 ne
rect 27154 30786 27246 30794
rect 27292 30827 27381 30832
tri 27381 30827 27389 30835 sw
rect 27292 30819 27389 30827
tri 27389 30819 27397 30827 sw
rect 27292 30811 27397 30819
tri 27397 30811 27405 30819 sw
rect 27292 30803 27405 30811
tri 27405 30803 27413 30811 sw
rect 70802 30804 71000 30862
rect 27292 30795 27413 30803
tri 27413 30795 27421 30803 sw
rect 27292 30787 27421 30795
tri 27421 30787 27429 30795 sw
rect 27292 30786 27429 30787
tri 27154 30778 27162 30786 ne
rect 27162 30783 27429 30786
tri 27429 30783 27433 30787 sw
rect 27162 30778 27433 30783
tri 27162 30770 27170 30778 ne
rect 27170 30775 27433 30778
tri 27433 30775 27441 30783 sw
rect 27170 30770 27441 30775
tri 27170 30768 27172 30770 ne
rect 27172 30768 27441 30770
tri 27172 30760 27180 30768 ne
rect 27180 30767 27441 30768
tri 27441 30767 27449 30775 sw
rect 27180 30760 27449 30767
tri 27180 30752 27188 30760 ne
rect 27188 30759 27449 30760
tri 27449 30759 27457 30767 sw
rect 27188 30752 27457 30759
tri 27188 30744 27196 30752 ne
rect 27196 30751 27457 30752
tri 27457 30751 27465 30759 sw
rect 70802 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
rect 27196 30744 27465 30751
tri 27196 30736 27204 30744 ne
rect 27204 30743 27465 30744
tri 27465 30743 27473 30751 sw
rect 27204 30736 27473 30743
tri 27204 30728 27212 30736 ne
rect 27212 30735 27473 30736
tri 27473 30735 27481 30743 sw
rect 27212 30728 27481 30735
tri 27212 30720 27220 30728 ne
rect 27220 30727 27481 30728
tri 27481 30727 27489 30735 sw
rect 27220 30720 27489 30727
tri 27220 30716 27224 30720 ne
rect 27224 30719 27489 30720
tri 27489 30719 27497 30727 sw
rect 27224 30716 27497 30719
tri 27497 30716 27500 30719 sw
tri 27224 30712 27228 30716 ne
rect 27228 30712 27500 30716
tri 27500 30712 27504 30716 sw
tri 27228 30704 27236 30712 ne
rect 27236 30711 27504 30712
tri 27504 30711 27505 30712 sw
rect 27236 30704 27505 30711
tri 27236 30696 27244 30704 ne
rect 27244 30703 27505 30704
tri 27505 30703 27513 30711 sw
rect 27244 30700 27513 30703
rect 27244 30696 27378 30700
tri 27244 30688 27252 30696 ne
rect 27252 30688 27378 30696
tri 27252 30680 27260 30688 ne
rect 27260 30680 27378 30688
tri 27260 30672 27268 30680 ne
rect 27268 30672 27378 30680
tri 27268 30664 27276 30672 ne
rect 27276 30664 27378 30672
tri 27276 30656 27284 30664 ne
rect 27284 30656 27378 30664
tri 27284 30648 27292 30656 ne
rect 27292 30654 27378 30656
rect 27424 30695 27513 30700
tri 27513 30695 27521 30703 sw
rect 70802 30700 71000 30758
rect 27424 30687 27521 30695
tri 27521 30687 27529 30695 sw
rect 27424 30679 27529 30687
tri 27529 30679 27537 30687 sw
rect 27424 30671 27537 30679
tri 27537 30671 27545 30679 sw
rect 27424 30663 27545 30671
tri 27545 30663 27553 30671 sw
rect 27424 30655 27553 30663
tri 27553 30655 27561 30663 sw
rect 27424 30654 27561 30655
rect 27292 30648 27561 30654
tri 27292 30640 27300 30648 ne
rect 27300 30647 27561 30648
tri 27561 30647 27569 30655 sw
rect 70802 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
rect 27300 30640 27569 30647
tri 27300 30632 27308 30640 ne
rect 27308 30639 27569 30640
tri 27569 30639 27577 30647 sw
rect 27308 30632 27577 30639
tri 27308 30624 27316 30632 ne
rect 27316 30631 27577 30632
tri 27577 30631 27585 30639 sw
rect 27316 30624 27585 30631
tri 27316 30616 27324 30624 ne
rect 27324 30623 27585 30624
tri 27585 30623 27593 30631 sw
rect 27324 30616 27593 30623
tri 27324 30608 27332 30616 ne
rect 27332 30615 27593 30616
tri 27593 30615 27601 30623 sw
rect 27332 30608 27601 30615
tri 27332 30600 27340 30608 ne
rect 27340 30607 27601 30608
tri 27601 30607 27609 30615 sw
rect 27340 30600 27609 30607
tri 27340 30592 27348 30600 ne
rect 27348 30599 27609 30600
tri 27609 30599 27617 30607 sw
rect 27348 30592 27617 30599
tri 27348 30584 27356 30592 ne
rect 27356 30591 27617 30592
tri 27617 30591 27625 30599 sw
rect 70802 30596 71000 30654
rect 27356 30584 27625 30591
tri 27356 30576 27364 30584 ne
rect 27364 30583 27625 30584
tri 27625 30583 27633 30591 sw
rect 27364 30576 27633 30583
tri 27633 30576 27640 30583 sw
tri 27364 30568 27372 30576 ne
rect 27372 30568 27640 30576
tri 27640 30568 27648 30576 sw
tri 27372 30560 27380 30568 ne
rect 27380 30560 27510 30568
tri 27380 30552 27388 30560 ne
rect 27388 30552 27510 30560
tri 27388 30544 27396 30552 ne
rect 27396 30544 27510 30552
tri 27396 30536 27404 30544 ne
rect 27404 30536 27510 30544
tri 27404 30528 27412 30536 ne
rect 27412 30528 27510 30536
tri 27412 30520 27420 30528 ne
rect 27420 30522 27510 30528
rect 27556 30560 27648 30568
tri 27648 30560 27656 30568 sw
rect 27556 30552 27656 30560
tri 27656 30552 27664 30560 sw
rect 27556 30544 27664 30552
tri 27664 30544 27672 30552 sw
rect 70802 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30536 27672 30544
tri 27672 30536 27680 30544 sw
rect 27556 30528 27680 30536
tri 27680 30528 27688 30536 sw
rect 27556 30522 27688 30528
rect 27420 30520 27688 30522
tri 27688 30520 27696 30528 sw
tri 27420 30512 27428 30520 ne
rect 27428 30512 27696 30520
tri 27696 30512 27704 30520 sw
tri 27428 30504 27436 30512 ne
rect 27436 30504 27704 30512
tri 27704 30504 27712 30512 sw
tri 27436 30496 27444 30504 ne
rect 27444 30496 27712 30504
tri 27712 30496 27720 30504 sw
tri 27444 30488 27452 30496 ne
rect 27452 30488 27720 30496
tri 27720 30488 27728 30496 sw
rect 70802 30492 71000 30550
tri 27452 30480 27460 30488 ne
rect 27460 30480 27728 30488
tri 27728 30480 27736 30488 sw
tri 27460 30472 27468 30480 ne
rect 27468 30472 27736 30480
tri 27736 30472 27744 30480 sw
tri 27468 30464 27476 30472 ne
rect 27476 30464 27744 30472
tri 27744 30464 27752 30472 sw
tri 27476 30456 27484 30464 ne
rect 27484 30456 27752 30464
tri 27752 30456 27760 30464 sw
tri 27484 30448 27492 30456 ne
rect 27492 30448 27760 30456
tri 27760 30448 27768 30456 sw
tri 27492 30440 27500 30448 ne
rect 27500 30440 27768 30448
tri 27768 30440 27776 30448 sw
rect 70802 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
tri 27500 30435 27505 30440 ne
rect 27505 30436 27776 30440
rect 27505 30435 27642 30436
tri 27505 30427 27513 30435 ne
rect 27513 30427 27642 30435
tri 27513 30419 27521 30427 ne
rect 27521 30419 27642 30427
tri 27521 30411 27529 30419 ne
rect 27529 30411 27642 30419
tri 27529 30403 27537 30411 ne
rect 27537 30403 27642 30411
tri 27537 30395 27545 30403 ne
rect 27545 30395 27642 30403
tri 27545 30387 27553 30395 ne
rect 27553 30390 27642 30395
rect 27688 30435 27776 30436
tri 27776 30435 27781 30440 sw
rect 27688 30427 27781 30435
tri 27781 30427 27789 30435 sw
rect 27688 30419 27789 30427
tri 27789 30419 27797 30427 sw
rect 27688 30411 27797 30419
tri 27797 30411 27805 30419 sw
rect 27688 30403 27805 30411
tri 27805 30403 27813 30411 sw
rect 27688 30395 27813 30403
tri 27813 30395 27821 30403 sw
rect 27688 30390 27821 30395
rect 27553 30387 27821 30390
tri 27821 30387 27829 30395 sw
rect 70802 30388 71000 30446
tri 27553 30379 27561 30387 ne
rect 27561 30379 27829 30387
tri 27829 30379 27837 30387 sw
tri 27561 30371 27569 30379 ne
rect 27569 30371 27837 30379
tri 27837 30371 27845 30379 sw
tri 27569 30363 27577 30371 ne
rect 27577 30363 27845 30371
tri 27845 30363 27853 30371 sw
tri 27577 30355 27585 30363 ne
rect 27585 30355 27853 30363
tri 27853 30355 27861 30363 sw
tri 27585 30347 27593 30355 ne
rect 27593 30347 27861 30355
tri 27861 30347 27869 30355 sw
tri 27593 30339 27601 30347 ne
rect 27601 30339 27869 30347
tri 27869 30339 27877 30347 sw
rect 70802 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27601 30331 27609 30339 ne
rect 27609 30331 27877 30339
tri 27877 30331 27885 30339 sw
tri 27609 30323 27617 30331 ne
rect 27617 30323 27885 30331
tri 27885 30323 27893 30331 sw
tri 27617 30315 27625 30323 ne
rect 27625 30315 27893 30323
tri 27893 30315 27901 30323 sw
tri 27625 30313 27627 30315 ne
rect 27627 30313 27901 30315
tri 27901 30313 27903 30315 sw
tri 27627 30305 27635 30313 ne
rect 27635 30305 27903 30313
tri 27903 30305 27911 30313 sw
tri 27635 30297 27643 30305 ne
rect 27643 30304 27911 30305
rect 27643 30297 27774 30304
tri 27643 30289 27651 30297 ne
rect 27651 30289 27774 30297
tri 27651 30281 27659 30289 ne
rect 27659 30281 27774 30289
tri 27659 30273 27667 30281 ne
rect 27667 30273 27774 30281
tri 27667 30265 27675 30273 ne
rect 27675 30265 27774 30273
tri 27675 30257 27683 30265 ne
rect 27683 30258 27774 30265
rect 27820 30297 27911 30304
tri 27911 30297 27919 30305 sw
rect 27820 30289 27919 30297
tri 27919 30289 27927 30297 sw
rect 27820 30281 27927 30289
tri 27927 30281 27935 30289 sw
rect 70802 30284 71000 30342
rect 27820 30273 27935 30281
tri 27935 30273 27943 30281 sw
rect 27820 30265 27943 30273
tri 27943 30265 27951 30273 sw
rect 27820 30258 27951 30265
rect 27683 30257 27951 30258
tri 27951 30257 27959 30265 sw
tri 27683 30249 27691 30257 ne
rect 27691 30249 27959 30257
tri 27959 30249 27967 30257 sw
tri 27691 30241 27699 30249 ne
rect 27699 30241 27967 30249
tri 27967 30241 27975 30249 sw
tri 27699 30233 27707 30241 ne
rect 27707 30233 27975 30241
tri 27975 30233 27983 30241 sw
rect 70802 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27707 30225 27715 30233 ne
rect 27715 30225 27983 30233
tri 27983 30225 27991 30233 sw
tri 27715 30217 27723 30225 ne
rect 27723 30217 27991 30225
tri 27991 30217 27999 30225 sw
tri 27723 30209 27731 30217 ne
rect 27731 30209 27999 30217
tri 27999 30209 28007 30217 sw
tri 27731 30207 27733 30209 ne
rect 27733 30207 28007 30209
tri 28007 30207 28009 30209 sw
tri 27733 30199 27741 30207 ne
rect 27741 30199 28009 30207
tri 28009 30199 28017 30207 sw
tri 27741 30191 27749 30199 ne
rect 27749 30191 28017 30199
tri 28017 30191 28025 30199 sw
tri 27749 30183 27757 30191 ne
rect 27757 30183 28025 30191
tri 28025 30183 28033 30191 sw
tri 27757 30175 27765 30183 ne
rect 27765 30175 28033 30183
tri 28033 30175 28041 30183 sw
rect 70802 30180 71000 30238
tri 27765 30167 27773 30175 ne
rect 27773 30172 28041 30175
rect 27773 30167 27906 30172
tri 27773 30159 27781 30167 ne
rect 27781 30159 27906 30167
tri 27781 30151 27789 30159 ne
rect 27789 30151 27906 30159
tri 27789 30143 27797 30151 ne
rect 27797 30143 27906 30151
tri 27797 30135 27805 30143 ne
rect 27805 30135 27906 30143
tri 27805 30127 27813 30135 ne
rect 27813 30127 27906 30135
tri 27813 30119 27821 30127 ne
rect 27821 30126 27906 30127
rect 27952 30167 28041 30172
tri 28041 30167 28049 30175 sw
rect 27952 30159 28049 30167
tri 28049 30159 28057 30167 sw
rect 27952 30151 28057 30159
tri 28057 30151 28065 30159 sw
rect 27952 30143 28065 30151
tri 28065 30143 28073 30151 sw
rect 27952 30135 28073 30143
tri 28073 30135 28081 30143 sw
rect 27952 30127 28081 30135
tri 28081 30127 28089 30135 sw
rect 70802 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 27952 30126 28089 30127
rect 27821 30119 28089 30126
tri 28089 30119 28097 30127 sw
tri 27821 30111 27829 30119 ne
rect 27829 30111 28097 30119
tri 28097 30111 28105 30119 sw
tri 27829 30103 27837 30111 ne
rect 27837 30103 28105 30111
tri 28105 30103 28113 30111 sw
tri 27837 30095 27845 30103 ne
rect 27845 30095 28113 30103
tri 28113 30095 28121 30103 sw
tri 27845 30087 27853 30095 ne
rect 27853 30087 28121 30095
tri 28121 30087 28129 30095 sw
tri 27853 30079 27861 30087 ne
rect 27861 30079 28129 30087
tri 28129 30079 28137 30087 sw
tri 27861 30071 27869 30079 ne
rect 27869 30071 28137 30079
tri 28137 30071 28145 30079 sw
rect 70802 30076 71000 30134
tri 27869 30063 27877 30071 ne
rect 27877 30063 28145 30071
tri 28145 30063 28153 30071 sw
tri 27877 30061 27879 30063 ne
rect 27879 30061 28153 30063
tri 28153 30061 28155 30063 sw
tri 27879 30053 27887 30061 ne
rect 27887 30053 28155 30061
tri 28155 30053 28163 30061 sw
tri 27887 30045 27895 30053 ne
rect 27895 30045 28163 30053
tri 28163 30045 28171 30053 sw
tri 27895 30037 27903 30045 ne
rect 27903 30040 28171 30045
rect 27903 30037 28038 30040
tri 27903 30029 27911 30037 ne
rect 27911 30029 28038 30037
tri 27911 30021 27919 30029 ne
rect 27919 30021 28038 30029
tri 27919 30013 27927 30021 ne
rect 27927 30013 28038 30021
tri 27927 30005 27935 30013 ne
rect 27935 30005 28038 30013
tri 27935 29997 27943 30005 ne
rect 27943 29997 28038 30005
tri 27943 29989 27951 29997 ne
rect 27951 29994 28038 29997
rect 28084 30037 28171 30040
tri 28171 30037 28179 30045 sw
rect 28084 30029 28179 30037
tri 28179 30029 28187 30037 sw
rect 70802 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 30021 28187 30029
tri 28187 30021 28195 30029 sw
rect 28084 30013 28195 30021
tri 28195 30013 28203 30021 sw
rect 28084 30005 28203 30013
tri 28203 30005 28211 30013 sw
rect 28084 29997 28211 30005
tri 28211 29997 28219 30005 sw
rect 28084 29994 28219 29997
rect 27951 29989 28219 29994
tri 28219 29989 28227 29997 sw
tri 27951 29981 27959 29989 ne
rect 27959 29981 28227 29989
tri 28227 29981 28235 29989 sw
tri 27959 29973 27967 29981 ne
rect 27967 29973 28235 29981
tri 28235 29973 28243 29981 sw
tri 27967 29965 27975 29973 ne
rect 27975 29965 28243 29973
tri 28243 29965 28251 29973 sw
rect 70802 29972 71000 30030
tri 27975 29957 27983 29965 ne
rect 27983 29957 28251 29965
tri 28251 29957 28259 29965 sw
tri 27983 29949 27991 29957 ne
rect 27991 29949 28259 29957
tri 28259 29949 28267 29957 sw
tri 27991 29941 27999 29949 ne
rect 27999 29941 28267 29949
tri 28267 29941 28275 29949 sw
tri 27999 29933 28007 29941 ne
rect 28007 29933 28275 29941
tri 28275 29933 28283 29941 sw
tri 28007 29925 28015 29933 ne
rect 28015 29925 28283 29933
tri 28283 29925 28291 29933 sw
rect 70802 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
tri 28015 29923 28017 29925 ne
rect 28017 29923 28291 29925
tri 28291 29923 28293 29925 sw
tri 28017 29915 28025 29923 ne
rect 28025 29915 28293 29923
tri 28293 29915 28301 29923 sw
tri 28025 29907 28033 29915 ne
rect 28033 29908 28301 29915
rect 28033 29907 28170 29908
tri 28033 29899 28041 29907 ne
rect 28041 29899 28170 29907
tri 28041 29891 28049 29899 ne
rect 28049 29891 28170 29899
tri 28049 29883 28057 29891 ne
rect 28057 29883 28170 29891
tri 28057 29875 28065 29883 ne
rect 28065 29875 28170 29883
tri 28065 29867 28073 29875 ne
rect 28073 29867 28170 29875
tri 28073 29859 28081 29867 ne
rect 28081 29862 28170 29867
rect 28216 29907 28301 29908
tri 28301 29907 28309 29915 sw
rect 28216 29899 28309 29907
tri 28309 29899 28317 29907 sw
rect 28216 29891 28317 29899
tri 28317 29891 28325 29899 sw
rect 28216 29883 28325 29891
tri 28325 29883 28333 29891 sw
rect 28216 29875 28333 29883
tri 28333 29875 28341 29883 sw
rect 28216 29867 28341 29875
tri 28341 29867 28349 29875 sw
rect 70802 29868 71000 29926
rect 28216 29862 28349 29867
rect 28081 29859 28349 29862
tri 28349 29859 28357 29867 sw
tri 28081 29851 28089 29859 ne
rect 28089 29851 28357 29859
tri 28357 29851 28365 29859 sw
tri 28089 29843 28097 29851 ne
rect 28097 29843 28365 29851
tri 28365 29843 28373 29851 sw
tri 28097 29835 28105 29843 ne
rect 28105 29835 28373 29843
tri 28373 29835 28381 29843 sw
tri 28105 29827 28113 29835 ne
rect 28113 29827 28381 29835
tri 28381 29827 28389 29835 sw
tri 28113 29819 28121 29827 ne
rect 28121 29819 28389 29827
tri 28389 29819 28397 29827 sw
rect 70802 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
tri 28121 29811 28129 29819 ne
rect 28129 29811 28397 29819
tri 28397 29811 28405 29819 sw
tri 28129 29803 28137 29811 ne
rect 28137 29803 28405 29811
tri 28405 29803 28413 29811 sw
tri 28137 29795 28145 29803 ne
rect 28145 29795 28413 29803
tri 28413 29795 28421 29803 sw
tri 28145 29787 28153 29795 ne
rect 28153 29787 28421 29795
tri 28421 29787 28429 29795 sw
tri 28153 29781 28159 29787 ne
rect 28159 29781 28429 29787
tri 28159 29773 28167 29781 ne
rect 28167 29780 28429 29781
tri 28429 29780 28436 29787 sw
rect 28167 29776 28436 29780
rect 28167 29773 28302 29776
tri 28167 29765 28175 29773 ne
rect 28175 29765 28302 29773
tri 28175 29757 28183 29765 ne
rect 28183 29757 28302 29765
tri 28183 29749 28191 29757 ne
rect 28191 29749 28302 29757
tri 28191 29741 28199 29749 ne
rect 28199 29741 28302 29749
tri 28199 29733 28207 29741 ne
rect 28207 29733 28302 29741
tri 28207 29725 28215 29733 ne
rect 28215 29730 28302 29733
rect 28348 29772 28436 29776
tri 28436 29772 28444 29780 sw
rect 28348 29764 28444 29772
tri 28444 29764 28452 29772 sw
rect 70802 29764 71000 29822
rect 28348 29756 28452 29764
tri 28452 29756 28460 29764 sw
rect 28348 29748 28460 29756
tri 28460 29748 28468 29756 sw
rect 28348 29740 28468 29748
tri 28468 29740 28476 29748 sw
rect 28348 29732 28476 29740
tri 28476 29732 28484 29740 sw
rect 28348 29730 28484 29732
rect 28215 29725 28484 29730
tri 28215 29717 28223 29725 ne
rect 28223 29724 28484 29725
tri 28484 29724 28492 29732 sw
rect 28223 29717 28492 29724
tri 28223 29709 28231 29717 ne
rect 28231 29716 28492 29717
tri 28492 29716 28500 29724 sw
rect 70802 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
rect 28231 29709 28500 29716
tri 28231 29701 28239 29709 ne
rect 28239 29708 28500 29709
tri 28500 29708 28508 29716 sw
rect 28239 29701 28508 29708
tri 28239 29693 28247 29701 ne
rect 28247 29700 28508 29701
tri 28508 29700 28516 29708 sw
rect 28247 29693 28516 29700
tri 28247 29685 28255 29693 ne
rect 28255 29692 28516 29693
tri 28516 29692 28524 29700 sw
rect 28255 29685 28524 29692
tri 28255 29677 28263 29685 ne
rect 28263 29684 28524 29685
tri 28524 29684 28532 29692 sw
rect 28263 29677 28532 29684
tri 28263 29669 28271 29677 ne
rect 28271 29676 28532 29677
tri 28532 29676 28540 29684 sw
rect 28271 29669 28540 29676
tri 28271 29661 28279 29669 ne
rect 28279 29668 28540 29669
tri 28540 29668 28548 29676 sw
rect 28279 29661 28548 29668
tri 28279 29657 28283 29661 ne
rect 28283 29660 28548 29661
tri 28548 29660 28556 29668 sw
rect 70802 29660 71000 29718
rect 28283 29657 28556 29660
tri 28556 29657 28559 29660 sw
tri 28283 29653 28287 29657 ne
rect 28287 29653 28559 29657
tri 28287 29645 28295 29653 ne
rect 28295 29652 28559 29653
tri 28559 29652 28564 29657 sw
rect 28295 29645 28564 29652
tri 28295 29637 28303 29645 ne
rect 28303 29644 28564 29645
tri 28564 29644 28572 29652 sw
rect 28303 29637 28434 29644
tri 28303 29629 28311 29637 ne
rect 28311 29629 28434 29637
tri 28311 29621 28319 29629 ne
rect 28319 29621 28434 29629
tri 28319 29613 28327 29621 ne
rect 28327 29613 28434 29621
tri 28327 29605 28335 29613 ne
rect 28335 29605 28434 29613
tri 28335 29597 28343 29605 ne
rect 28343 29598 28434 29605
rect 28480 29636 28572 29644
tri 28572 29636 28580 29644 sw
rect 28480 29628 28580 29636
tri 28580 29628 28588 29636 sw
rect 28480 29620 28588 29628
tri 28588 29620 28596 29628 sw
rect 28480 29612 28596 29620
tri 28596 29612 28604 29620 sw
rect 70802 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 28480 29604 28604 29612
tri 28604 29604 28612 29612 sw
rect 28480 29598 28612 29604
rect 28343 29597 28612 29598
tri 28343 29589 28351 29597 ne
rect 28351 29596 28612 29597
tri 28612 29596 28620 29604 sw
rect 28351 29589 28620 29596
tri 28351 29581 28359 29589 ne
rect 28359 29588 28620 29589
tri 28620 29588 28628 29596 sw
rect 28359 29581 28628 29588
tri 28359 29573 28367 29581 ne
rect 28367 29580 28628 29581
tri 28628 29580 28636 29588 sw
rect 28367 29573 28636 29580
tri 28367 29565 28375 29573 ne
rect 28375 29572 28636 29573
tri 28636 29572 28644 29580 sw
rect 28375 29565 28644 29572
tri 28375 29557 28383 29565 ne
rect 28383 29564 28644 29565
tri 28644 29564 28652 29572 sw
rect 28383 29557 28652 29564
tri 28383 29549 28391 29557 ne
rect 28391 29556 28652 29557
tri 28652 29556 28660 29564 sw
rect 70802 29556 71000 29614
rect 28391 29549 28660 29556
tri 28391 29541 28399 29549 ne
rect 28399 29548 28660 29549
tri 28660 29548 28668 29556 sw
rect 28399 29541 28668 29548
tri 28399 29533 28407 29541 ne
rect 28407 29540 28668 29541
tri 28668 29540 28676 29548 sw
rect 28407 29533 28676 29540
tri 28407 29525 28415 29533 ne
rect 28415 29532 28676 29533
tri 28676 29532 28684 29540 sw
rect 28415 29525 28684 29532
tri 28415 29517 28423 29525 ne
rect 28423 29524 28684 29525
tri 28684 29524 28692 29532 sw
rect 28423 29521 28692 29524
tri 28692 29521 28695 29524 sw
rect 28423 29517 28695 29521
tri 28423 29513 28427 29517 ne
rect 28427 29513 28695 29517
tri 28695 29513 28703 29521 sw
tri 28427 29505 28435 29513 ne
rect 28435 29512 28703 29513
rect 28435 29505 28566 29512
tri 28435 29497 28443 29505 ne
rect 28443 29497 28566 29505
tri 28443 29489 28451 29497 ne
rect 28451 29489 28566 29497
tri 28451 29481 28459 29489 ne
rect 28459 29481 28566 29489
tri 28459 29473 28467 29481 ne
rect 28467 29473 28566 29481
tri 28467 29465 28475 29473 ne
rect 28475 29466 28566 29473
rect 28612 29505 28703 29512
tri 28703 29505 28711 29513 sw
rect 70802 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29497 28711 29505
tri 28711 29497 28719 29505 sw
rect 28612 29489 28719 29497
tri 28719 29489 28727 29497 sw
rect 28612 29481 28727 29489
tri 28727 29481 28735 29489 sw
rect 28612 29473 28735 29481
tri 28735 29473 28743 29481 sw
rect 28612 29466 28743 29473
rect 28475 29465 28743 29466
tri 28743 29465 28751 29473 sw
tri 28475 29457 28483 29465 ne
rect 28483 29457 28751 29465
tri 28751 29457 28759 29465 sw
tri 28483 29449 28491 29457 ne
rect 28491 29449 28759 29457
tri 28759 29449 28767 29457 sw
rect 70802 29452 71000 29510
tri 28491 29441 28499 29449 ne
rect 28499 29441 28767 29449
tri 28767 29441 28775 29449 sw
tri 28499 29433 28507 29441 ne
rect 28507 29433 28775 29441
tri 28775 29433 28783 29441 sw
tri 28507 29425 28515 29433 ne
rect 28515 29425 28783 29433
tri 28783 29425 28791 29433 sw
tri 28515 29417 28523 29425 ne
rect 28523 29417 28791 29425
tri 28791 29417 28799 29425 sw
tri 28523 29409 28531 29417 ne
rect 28531 29409 28799 29417
tri 28799 29409 28807 29417 sw
tri 28531 29401 28539 29409 ne
rect 28539 29401 28807 29409
tri 28807 29401 28815 29409 sw
rect 70802 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28539 29393 28547 29401 ne
rect 28547 29393 28815 29401
tri 28815 29393 28823 29401 sw
tri 28547 29385 28555 29393 ne
rect 28555 29385 28823 29393
tri 28823 29385 28831 29393 sw
tri 28555 29381 28559 29385 ne
rect 28559 29381 28831 29385
tri 28831 29381 28835 29385 sw
tri 28559 29377 28563 29381 ne
rect 28563 29380 28835 29381
rect 28563 29377 28698 29380
tri 28563 29369 28571 29377 ne
rect 28571 29369 28698 29377
tri 28571 29361 28579 29369 ne
rect 28579 29361 28698 29369
tri 28579 29353 28587 29361 ne
rect 28587 29353 28698 29361
tri 28587 29345 28595 29353 ne
rect 28595 29345 28698 29353
tri 28595 29337 28603 29345 ne
rect 28603 29337 28698 29345
tri 28603 29329 28611 29337 ne
rect 28611 29334 28698 29337
rect 28744 29377 28835 29380
tri 28835 29377 28839 29381 sw
rect 28744 29369 28839 29377
tri 28839 29369 28847 29377 sw
rect 28744 29361 28847 29369
tri 28847 29361 28855 29369 sw
rect 28744 29353 28855 29361
tri 28855 29353 28863 29361 sw
rect 28744 29345 28863 29353
tri 28863 29345 28871 29353 sw
rect 70802 29348 71000 29406
rect 28744 29337 28871 29345
tri 28871 29337 28879 29345 sw
rect 28744 29334 28879 29337
rect 28611 29329 28879 29334
tri 28879 29329 28887 29337 sw
tri 28611 29321 28619 29329 ne
rect 28619 29321 28887 29329
tri 28887 29321 28895 29329 sw
tri 28619 29313 28627 29321 ne
rect 28627 29313 28895 29321
tri 28895 29313 28903 29321 sw
tri 28627 29305 28635 29313 ne
rect 28635 29305 28903 29313
tri 28903 29305 28911 29313 sw
tri 28635 29297 28643 29305 ne
rect 28643 29297 28911 29305
tri 28911 29297 28919 29305 sw
rect 70802 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28643 29289 28651 29297 ne
rect 28651 29289 28919 29297
tri 28919 29289 28927 29297 sw
tri 28651 29281 28659 29289 ne
rect 28659 29281 28927 29289
tri 28927 29281 28935 29289 sw
tri 28659 29273 28667 29281 ne
rect 28667 29273 28935 29281
tri 28935 29273 28943 29281 sw
tri 28667 29265 28675 29273 ne
rect 28675 29265 28943 29273
tri 28943 29265 28951 29273 sw
tri 28675 29257 28683 29265 ne
rect 28683 29257 28951 29265
tri 28951 29257 28959 29265 sw
tri 28683 29249 28691 29257 ne
rect 28691 29256 28959 29257
tri 28959 29256 28960 29257 sw
rect 28691 29249 28960 29256
tri 28691 29242 28698 29249 ne
rect 28698 29248 28960 29249
tri 28960 29248 28968 29256 sw
rect 28698 29242 28830 29248
tri 28698 29234 28706 29242 ne
rect 28706 29234 28830 29242
tri 28706 29226 28714 29234 ne
rect 28714 29226 28830 29234
tri 28714 29218 28722 29226 ne
rect 28722 29218 28830 29226
tri 28722 29210 28730 29218 ne
rect 28730 29210 28830 29218
tri 28730 29202 28738 29210 ne
rect 28738 29202 28830 29210
rect 28876 29240 28968 29248
tri 28968 29240 28976 29248 sw
rect 70802 29244 71000 29302
rect 28876 29232 28976 29240
tri 28976 29232 28984 29240 sw
rect 28876 29224 28984 29232
tri 28984 29224 28992 29232 sw
rect 28876 29216 28992 29224
tri 28992 29216 29000 29224 sw
rect 28876 29208 29000 29216
tri 29000 29208 29008 29216 sw
rect 28876 29202 29008 29208
tri 28738 29194 28746 29202 ne
rect 28746 29200 29008 29202
tri 29008 29200 29016 29208 sw
rect 28746 29194 29016 29200
tri 28746 29186 28754 29194 ne
rect 28754 29192 29016 29194
tri 29016 29192 29024 29200 sw
rect 70802 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
rect 28754 29186 29024 29192
tri 28754 29178 28762 29186 ne
rect 28762 29184 29024 29186
tri 29024 29184 29032 29192 sw
rect 28762 29178 29032 29184
tri 28762 29170 28770 29178 ne
rect 28770 29176 29032 29178
tri 29032 29176 29040 29184 sw
rect 28770 29170 29040 29176
tri 28770 29162 28778 29170 ne
rect 28778 29168 29040 29170
tri 29040 29168 29048 29176 sw
rect 28778 29162 29048 29168
tri 28778 29154 28786 29162 ne
rect 28786 29160 29048 29162
tri 29048 29160 29056 29168 sw
rect 28786 29154 29056 29160
tri 28786 29146 28794 29154 ne
rect 28794 29152 29056 29154
tri 29056 29152 29064 29160 sw
rect 28794 29146 29064 29152
tri 28794 29138 28802 29146 ne
rect 28802 29144 29064 29146
tri 29064 29144 29072 29152 sw
rect 28802 29138 29072 29144
tri 28802 29130 28810 29138 ne
rect 28810 29136 29072 29138
tri 29072 29136 29080 29144 sw
rect 70802 29140 71000 29198
rect 28810 29130 29080 29136
tri 28810 29122 28818 29130 ne
rect 28818 29128 29080 29130
tri 29080 29128 29088 29136 sw
rect 28818 29124 29088 29128
tri 29088 29124 29092 29128 sw
rect 28818 29122 29092 29124
tri 28818 29114 28826 29122 ne
rect 28826 29120 29092 29122
tri 29092 29120 29096 29124 sw
rect 28826 29116 29096 29120
rect 28826 29114 28962 29116
tri 28826 29110 28830 29114 ne
rect 28830 29110 28962 29114
tri 28830 29106 28834 29110 ne
rect 28834 29106 28962 29110
tri 28834 29098 28842 29106 ne
rect 28842 29098 28962 29106
tri 28842 29090 28850 29098 ne
rect 28850 29090 28962 29098
tri 28850 29082 28858 29090 ne
rect 28858 29082 28962 29090
tri 28858 29074 28866 29082 ne
rect 28866 29074 28962 29082
tri 28866 29066 28874 29074 ne
rect 28874 29070 28962 29074
rect 29008 29112 29096 29116
tri 29096 29112 29104 29120 sw
rect 29008 29104 29104 29112
tri 29104 29104 29112 29112 sw
rect 29008 29096 29112 29104
tri 29112 29096 29120 29104 sw
rect 29008 29088 29120 29096
tri 29120 29088 29128 29096 sw
rect 70802 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 29008 29080 29128 29088
tri 29128 29080 29136 29088 sw
rect 29008 29072 29136 29080
tri 29136 29072 29144 29080 sw
rect 29008 29071 29144 29072
tri 29144 29071 29145 29072 sw
rect 29008 29070 29145 29071
rect 28874 29066 29145 29070
tri 28874 29058 28882 29066 ne
rect 28882 29063 29145 29066
tri 29145 29063 29153 29071 sw
rect 28882 29058 29153 29063
tri 28882 29057 28883 29058 ne
rect 28883 29057 29153 29058
tri 28883 29049 28891 29057 ne
rect 28891 29055 29153 29057
tri 29153 29055 29161 29063 sw
rect 28891 29049 29161 29055
tri 28891 29041 28899 29049 ne
rect 28899 29047 29161 29049
tri 29161 29047 29169 29055 sw
rect 28899 29041 29169 29047
tri 28899 29033 28907 29041 ne
rect 28907 29039 29169 29041
tri 29169 29039 29177 29047 sw
rect 28907 29033 29177 29039
tri 28907 29025 28915 29033 ne
rect 28915 29031 29177 29033
tri 29177 29031 29185 29039 sw
rect 70802 29036 71000 29094
rect 28915 29025 29185 29031
tri 28915 29017 28923 29025 ne
rect 28923 29023 29185 29025
tri 29185 29023 29193 29031 sw
rect 28923 29017 29193 29023
tri 28923 29009 28931 29017 ne
rect 28931 29015 29193 29017
tri 29193 29015 29201 29023 sw
rect 28931 29009 29201 29015
tri 28931 29001 28939 29009 ne
rect 28939 29007 29201 29009
tri 29201 29007 29209 29015 sw
rect 28939 29001 29209 29007
tri 28939 28993 28947 29001 ne
rect 28947 28999 29209 29001
tri 29209 28999 29217 29007 sw
rect 28947 28993 29217 28999
tri 28947 28985 28955 28993 ne
rect 28955 28991 29217 28993
tri 29217 28991 29225 28999 sw
rect 28955 28985 29225 28991
tri 28955 28977 28963 28985 ne
rect 28963 28984 29225 28985
rect 28963 28977 29094 28984
tri 28963 28969 28971 28977 ne
rect 28971 28969 29094 28977
tri 28971 28961 28979 28969 ne
rect 28979 28961 29094 28969
tri 28979 28953 28987 28961 ne
rect 28987 28953 29094 28961
tri 28987 28945 28995 28953 ne
rect 28995 28945 29094 28953
tri 28995 28937 29003 28945 ne
rect 29003 28938 29094 28945
rect 29140 28983 29225 28984
tri 29225 28983 29233 28991 sw
rect 70802 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 29140 28975 29233 28983
tri 29233 28975 29241 28983 sw
rect 29140 28967 29241 28975
tri 29241 28967 29249 28975 sw
rect 29140 28959 29249 28967
tri 29249 28959 29257 28967 sw
rect 29140 28951 29257 28959
tri 29257 28951 29265 28959 sw
rect 29140 28946 29265 28951
tri 29265 28946 29270 28951 sw
rect 29140 28938 29270 28946
tri 29270 28938 29278 28946 sw
rect 29003 28937 29278 28938
tri 29003 28929 29011 28937 ne
rect 29011 28930 29278 28937
tri 29278 28930 29286 28938 sw
rect 70802 28932 71000 28990
rect 29011 28929 29286 28930
tri 29011 28922 29018 28929 ne
rect 29018 28922 29286 28929
tri 29286 28922 29294 28930 sw
tri 29018 28914 29026 28922 ne
rect 29026 28914 29294 28922
tri 29294 28914 29302 28922 sw
tri 29026 28906 29034 28914 ne
rect 29034 28906 29302 28914
tri 29302 28906 29310 28914 sw
tri 29034 28898 29042 28906 ne
rect 29042 28898 29310 28906
tri 29310 28898 29318 28906 sw
tri 29042 28890 29050 28898 ne
rect 29050 28890 29318 28898
tri 29318 28890 29326 28898 sw
tri 29050 28882 29058 28890 ne
rect 29058 28882 29326 28890
tri 29326 28882 29334 28890 sw
rect 70802 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29058 28874 29066 28882 ne
rect 29066 28874 29334 28882
tri 29334 28874 29342 28882 sw
tri 29066 28866 29074 28874 ne
rect 29074 28866 29342 28874
tri 29342 28866 29350 28874 sw
tri 29074 28858 29082 28866 ne
rect 29082 28863 29350 28866
tri 29350 28863 29353 28866 sw
rect 29082 28858 29353 28863
tri 29082 28850 29090 28858 ne
rect 29090 28855 29353 28858
tri 29353 28855 29361 28863 sw
rect 29090 28852 29361 28855
rect 29090 28850 29226 28852
tri 29090 28846 29094 28850 ne
rect 29094 28846 29226 28850
tri 29094 28842 29098 28846 ne
rect 29098 28842 29226 28846
tri 29098 28834 29106 28842 ne
rect 29106 28834 29226 28842
tri 29106 28826 29114 28834 ne
rect 29114 28826 29226 28834
tri 29114 28818 29122 28826 ne
rect 29122 28818 29226 28826
tri 29122 28810 29130 28818 ne
rect 29130 28810 29226 28818
tri 29130 28802 29138 28810 ne
rect 29138 28806 29226 28810
rect 29272 28847 29361 28852
tri 29361 28847 29369 28855 sw
rect 29272 28842 29369 28847
tri 29369 28842 29374 28847 sw
rect 29272 28839 29374 28842
tri 29374 28839 29377 28842 sw
rect 29272 28831 29377 28839
tri 29377 28831 29385 28839 sw
rect 29272 28823 29385 28831
tri 29385 28823 29393 28831 sw
rect 70802 28828 71000 28886
rect 29272 28815 29393 28823
tri 29393 28815 29401 28823 sw
rect 29272 28807 29401 28815
tri 29401 28807 29409 28815 sw
rect 29272 28806 29409 28807
rect 29138 28802 29409 28806
tri 29138 28794 29146 28802 ne
rect 29146 28799 29409 28802
tri 29409 28799 29417 28807 sw
rect 29146 28798 29417 28799
tri 29417 28798 29418 28799 sw
rect 29146 28794 29418 28798
tri 29146 28786 29154 28794 ne
rect 29154 28790 29418 28794
tri 29418 28790 29426 28798 sw
rect 29154 28786 29426 28790
tri 29154 28783 29157 28786 ne
rect 29157 28783 29426 28786
tri 29157 28775 29165 28783 ne
rect 29165 28782 29426 28783
tri 29426 28782 29434 28790 sw
rect 70802 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 29165 28775 29434 28782
tri 29165 28767 29173 28775 ne
rect 29173 28774 29434 28775
tri 29434 28774 29442 28782 sw
rect 29173 28767 29442 28774
tri 29173 28759 29181 28767 ne
rect 29181 28766 29442 28767
tri 29442 28766 29450 28774 sw
rect 29181 28759 29450 28766
tri 29181 28751 29189 28759 ne
rect 29189 28758 29450 28759
tri 29450 28758 29458 28766 sw
rect 29189 28751 29458 28758
tri 29189 28743 29197 28751 ne
rect 29197 28750 29458 28751
tri 29458 28750 29466 28758 sw
rect 29197 28743 29466 28750
tri 29197 28735 29205 28743 ne
rect 29205 28742 29466 28743
tri 29466 28742 29474 28750 sw
rect 29205 28735 29474 28742
tri 29205 28727 29213 28735 ne
rect 29213 28734 29474 28735
tri 29474 28734 29482 28742 sw
rect 29213 28727 29482 28734
tri 29213 28719 29221 28727 ne
rect 29221 28726 29482 28727
tri 29482 28726 29490 28734 sw
rect 29221 28720 29490 28726
rect 29221 28719 29358 28720
tri 29221 28711 29229 28719 ne
rect 29229 28711 29358 28719
tri 29229 28703 29237 28711 ne
rect 29237 28703 29358 28711
tri 29237 28695 29245 28703 ne
rect 29245 28695 29358 28703
tri 29245 28687 29253 28695 ne
rect 29253 28687 29358 28695
tri 29253 28679 29261 28687 ne
rect 29261 28679 29358 28687
tri 29261 28671 29269 28679 ne
rect 29269 28674 29358 28679
rect 29404 28718 29490 28720
tri 29490 28718 29498 28726 sw
rect 70802 28724 71000 28782
rect 29404 28710 29498 28718
tri 29498 28710 29506 28718 sw
rect 29404 28702 29506 28710
tri 29506 28702 29514 28710 sw
rect 29404 28694 29514 28702
tri 29514 28694 29522 28702 sw
rect 29404 28686 29522 28694
tri 29522 28686 29530 28694 sw
rect 29404 28678 29530 28686
tri 29530 28678 29538 28686 sw
rect 70802 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 29404 28674 29538 28678
rect 29269 28671 29538 28674
tri 29269 28663 29277 28671 ne
rect 29277 28670 29538 28671
tri 29538 28670 29546 28678 sw
rect 29277 28663 29546 28670
tri 29277 28655 29285 28663 ne
rect 29285 28662 29546 28663
tri 29546 28662 29554 28670 sw
rect 29285 28655 29554 28662
tri 29285 28654 29286 28655 ne
rect 29286 28654 29554 28655
tri 29554 28654 29562 28662 sw
tri 29286 28646 29294 28654 ne
rect 29294 28646 29562 28654
tri 29562 28646 29570 28654 sw
tri 29294 28638 29302 28646 ne
rect 29302 28638 29570 28646
tri 29570 28638 29578 28646 sw
tri 29302 28630 29310 28638 ne
rect 29310 28630 29578 28638
tri 29578 28630 29586 28638 sw
tri 29310 28622 29318 28630 ne
rect 29318 28622 29586 28630
tri 29586 28622 29594 28630 sw
tri 29318 28614 29326 28622 ne
rect 29326 28614 29594 28622
tri 29594 28614 29602 28622 sw
rect 70802 28620 71000 28678
tri 29326 28606 29334 28614 ne
rect 29334 28606 29602 28614
tri 29602 28606 29610 28614 sw
tri 29334 28598 29342 28606 ne
rect 29342 28598 29610 28606
tri 29610 28598 29618 28606 sw
tri 29342 28590 29350 28598 ne
rect 29350 28590 29618 28598
tri 29618 28590 29626 28598 sw
tri 29350 28582 29358 28590 ne
rect 29358 28588 29626 28590
rect 29358 28582 29490 28588
tri 29358 28574 29366 28582 ne
rect 29366 28574 29490 28582
tri 29366 28571 29369 28574 ne
rect 29369 28571 29490 28574
tri 29369 28563 29377 28571 ne
rect 29377 28563 29490 28571
tri 29377 28555 29385 28563 ne
rect 29385 28555 29490 28563
tri 29385 28547 29393 28555 ne
rect 29393 28547 29490 28555
tri 29393 28539 29401 28547 ne
rect 29401 28542 29490 28547
rect 29536 28582 29626 28588
tri 29626 28582 29634 28590 sw
rect 29536 28579 29634 28582
tri 29634 28579 29637 28582 sw
rect 29536 28571 29637 28579
tri 29637 28571 29645 28579 sw
rect 70802 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28563 29645 28571
tri 29645 28563 29653 28571 sw
rect 29536 28555 29653 28563
tri 29653 28555 29661 28563 sw
rect 29536 28547 29661 28555
tri 29661 28547 29669 28555 sw
rect 29536 28542 29669 28547
rect 29401 28539 29669 28542
tri 29669 28539 29677 28547 sw
tri 29401 28531 29409 28539 ne
rect 29409 28531 29677 28539
tri 29677 28531 29685 28539 sw
tri 29409 28523 29417 28531 ne
rect 29417 28523 29685 28531
tri 29685 28523 29693 28531 sw
tri 29417 28515 29425 28523 ne
rect 29425 28515 29693 28523
tri 29693 28515 29701 28523 sw
rect 70802 28516 71000 28574
tri 29425 28507 29433 28515 ne
rect 29433 28514 29701 28515
tri 29701 28514 29702 28515 sw
rect 29433 28507 29702 28514
tri 29433 28503 29437 28507 ne
rect 29437 28506 29702 28507
tri 29702 28506 29710 28514 sw
rect 29437 28503 29710 28506
tri 29437 28495 29445 28503 ne
rect 29445 28498 29710 28503
tri 29710 28498 29718 28506 sw
rect 29445 28495 29718 28498
tri 29445 28487 29453 28495 ne
rect 29453 28490 29718 28495
tri 29718 28490 29726 28498 sw
rect 29453 28487 29726 28490
tri 29453 28479 29461 28487 ne
rect 29461 28482 29726 28487
tri 29726 28482 29734 28490 sw
rect 29461 28479 29734 28482
tri 29461 28471 29469 28479 ne
rect 29469 28474 29734 28479
tri 29734 28474 29742 28482 sw
rect 29469 28471 29742 28474
tri 29469 28463 29477 28471 ne
rect 29477 28466 29742 28471
tri 29742 28466 29750 28474 sw
rect 70802 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29477 28463 29750 28466
tri 29477 28455 29485 28463 ne
rect 29485 28458 29750 28463
tri 29750 28458 29758 28466 sw
rect 29485 28456 29758 28458
rect 29485 28455 29622 28456
tri 29485 28447 29493 28455 ne
rect 29493 28447 29622 28455
tri 29493 28439 29501 28447 ne
rect 29501 28439 29622 28447
tri 29501 28431 29509 28439 ne
rect 29509 28431 29622 28439
tri 29509 28423 29517 28431 ne
rect 29517 28423 29622 28431
tri 29517 28415 29525 28423 ne
rect 29525 28415 29622 28423
tri 29525 28407 29533 28415 ne
rect 29533 28410 29622 28415
rect 29668 28450 29758 28456
tri 29758 28450 29766 28458 sw
rect 29668 28442 29766 28450
tri 29766 28442 29774 28450 sw
rect 29668 28434 29774 28442
tri 29774 28434 29782 28442 sw
rect 29668 28426 29782 28434
tri 29782 28426 29790 28434 sw
rect 29668 28418 29790 28426
tri 29790 28418 29798 28426 sw
rect 29668 28411 29798 28418
tri 29798 28411 29805 28418 sw
rect 70802 28412 71000 28470
rect 29668 28410 29805 28411
rect 29533 28407 29805 28410
tri 29533 28399 29541 28407 ne
rect 29541 28403 29805 28407
tri 29805 28403 29813 28411 sw
rect 29541 28399 29813 28403
tri 29541 28391 29549 28399 ne
rect 29549 28395 29813 28399
tri 29813 28395 29821 28403 sw
rect 29549 28391 29821 28395
tri 29549 28386 29554 28391 ne
rect 29554 28387 29821 28391
tri 29821 28387 29829 28395 sw
rect 29554 28386 29829 28387
tri 29554 28378 29562 28386 ne
rect 29562 28379 29829 28386
tri 29829 28379 29837 28387 sw
rect 29562 28378 29837 28379
tri 29562 28370 29570 28378 ne
rect 29570 28371 29837 28378
tri 29837 28371 29845 28379 sw
rect 29570 28370 29845 28371
tri 29570 28362 29578 28370 ne
rect 29578 28363 29845 28370
tri 29845 28363 29853 28371 sw
rect 70802 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
rect 29578 28362 29853 28363
tri 29578 28354 29586 28362 ne
rect 29586 28355 29853 28362
tri 29853 28355 29861 28363 sw
rect 29586 28354 29861 28355
tri 29586 28346 29594 28354 ne
rect 29594 28347 29861 28354
tri 29861 28347 29869 28355 sw
rect 29594 28346 29869 28347
tri 29594 28338 29602 28346 ne
rect 29602 28339 29869 28346
tri 29869 28339 29877 28347 sw
rect 29602 28338 29877 28339
tri 29602 28330 29610 28338 ne
rect 29610 28335 29877 28338
tri 29877 28335 29881 28339 sw
rect 29610 28330 29881 28335
tri 29610 28322 29618 28330 ne
rect 29618 28327 29881 28330
tri 29881 28327 29889 28335 sw
rect 29618 28324 29889 28327
rect 29618 28322 29754 28324
tri 29618 28318 29622 28322 ne
rect 29622 28318 29754 28322
tri 29622 28314 29626 28318 ne
rect 29626 28314 29754 28318
tri 29626 28306 29634 28314 ne
rect 29634 28306 29754 28314
tri 29634 28298 29642 28306 ne
rect 29642 28298 29754 28306
tri 29642 28290 29650 28298 ne
rect 29650 28290 29754 28298
tri 29650 28282 29658 28290 ne
rect 29658 28282 29754 28290
tri 29658 28274 29666 28282 ne
rect 29666 28278 29754 28282
rect 29800 28319 29889 28324
tri 29889 28319 29897 28327 sw
rect 29800 28314 29897 28319
tri 29897 28314 29902 28319 sw
rect 29800 28306 29902 28314
tri 29902 28306 29910 28314 sw
rect 70802 28308 71000 28366
rect 29800 28298 29910 28306
tri 29910 28298 29918 28306 sw
rect 29800 28290 29918 28298
tri 29918 28290 29926 28298 sw
rect 29800 28282 29926 28290
tri 29926 28282 29934 28290 sw
rect 29800 28278 29934 28282
rect 29666 28274 29934 28278
tri 29934 28274 29942 28282 sw
tri 29666 28266 29674 28274 ne
rect 29674 28272 29942 28274
tri 29942 28272 29944 28274 sw
rect 29674 28266 29944 28272
tri 29674 28258 29682 28266 ne
rect 29682 28264 29944 28266
tri 29944 28264 29952 28272 sw
rect 29682 28258 29952 28264
tri 29682 28250 29690 28258 ne
rect 29690 28256 29952 28258
tri 29952 28256 29960 28264 sw
rect 70802 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
rect 29690 28250 29960 28256
tri 29690 28243 29697 28250 ne
rect 29697 28248 29960 28250
tri 29960 28248 29968 28256 sw
rect 29697 28243 29968 28248
tri 29697 28235 29705 28243 ne
rect 29705 28240 29968 28243
tri 29968 28240 29976 28248 sw
rect 29705 28235 29976 28240
tri 29705 28227 29713 28235 ne
rect 29713 28232 29976 28235
tri 29976 28232 29984 28240 sw
rect 29713 28227 29984 28232
tri 29713 28219 29721 28227 ne
rect 29721 28224 29984 28227
tri 29984 28224 29992 28232 sw
rect 29721 28219 29992 28224
tri 29721 28211 29729 28219 ne
rect 29729 28216 29992 28219
tri 29992 28216 30000 28224 sw
rect 29729 28211 30000 28216
tri 29729 28203 29737 28211 ne
rect 29737 28208 30000 28211
tri 30000 28208 30008 28216 sw
rect 29737 28203 30008 28208
tri 29737 28195 29745 28203 ne
rect 29745 28200 30008 28203
tri 30008 28200 30016 28208 sw
rect 70802 28204 71000 28262
rect 29745 28195 30016 28200
tri 29745 28187 29753 28195 ne
rect 29753 28192 30016 28195
tri 30016 28192 30024 28200 sw
rect 29753 28187 29886 28192
tri 29753 28179 29761 28187 ne
rect 29761 28179 29886 28187
tri 29761 28171 29769 28179 ne
rect 29769 28171 29886 28179
tri 29769 28163 29777 28171 ne
rect 29777 28163 29886 28171
tri 29777 28155 29785 28163 ne
rect 29785 28155 29886 28163
tri 29785 28147 29793 28155 ne
rect 29793 28147 29886 28155
tri 29793 28139 29801 28147 ne
rect 29801 28146 29886 28147
rect 29932 28184 30024 28192
tri 30024 28184 30032 28192 sw
rect 29932 28176 30032 28184
tri 30032 28176 30040 28184 sw
rect 29932 28168 30040 28176
tri 30040 28168 30048 28176 sw
rect 29932 28160 30048 28168
tri 30048 28160 30056 28168 sw
rect 29932 28152 30056 28160
tri 30056 28152 30064 28160 sw
rect 70802 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 29932 28151 30064 28152
tri 30064 28151 30065 28152 sw
rect 29932 28146 30065 28151
rect 29801 28143 30065 28146
tri 30065 28143 30073 28151 sw
rect 29801 28139 30073 28143
tri 29801 28131 29809 28139 ne
rect 29809 28135 30073 28139
tri 30073 28135 30081 28143 sw
rect 29809 28131 30081 28135
tri 29809 28123 29817 28131 ne
rect 29817 28127 30081 28131
tri 30081 28127 30089 28135 sw
rect 29817 28123 30089 28127
tri 29817 28115 29825 28123 ne
rect 29825 28119 30089 28123
tri 30089 28119 30097 28127 sw
rect 29825 28115 30097 28119
tri 29825 28107 29833 28115 ne
rect 29833 28111 30097 28115
tri 30097 28111 30105 28119 sw
rect 29833 28107 30105 28111
tri 29833 28099 29841 28107 ne
rect 29841 28103 30105 28107
tri 30105 28103 30113 28111 sw
rect 29841 28099 30113 28103
tri 29841 28091 29849 28099 ne
rect 29849 28095 30113 28099
tri 30113 28095 30121 28103 sw
rect 70802 28100 71000 28158
rect 29849 28091 30121 28095
tri 29849 28083 29857 28091 ne
rect 29857 28087 30121 28091
tri 30121 28087 30129 28095 sw
rect 29857 28083 30129 28087
tri 29857 28075 29865 28083 ne
rect 29865 28079 30129 28083
tri 30129 28079 30137 28087 sw
rect 29865 28075 30137 28079
tri 29865 28067 29873 28075 ne
rect 29873 28071 30137 28075
tri 30137 28071 30145 28079 sw
rect 29873 28067 30145 28071
tri 29873 28059 29881 28067 ne
rect 29881 28063 30145 28067
tri 30145 28063 30153 28071 sw
rect 29881 28060 30153 28063
rect 29881 28059 30018 28060
tri 29881 28051 29889 28059 ne
rect 29889 28051 30018 28059
tri 29889 28043 29897 28051 ne
rect 29897 28043 30018 28051
tri 29897 28035 29905 28043 ne
rect 29905 28035 30018 28043
tri 29905 28027 29913 28035 ne
rect 29913 28027 30018 28035
tri 29913 28019 29921 28027 ne
rect 29921 28019 30018 28027
tri 29921 28011 29929 28019 ne
rect 29929 28014 30018 28019
rect 30064 28055 30153 28060
tri 30153 28055 30161 28063 sw
rect 30064 28051 30161 28055
tri 30161 28051 30165 28055 sw
rect 70802 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28043 30165 28051
tri 30165 28043 30173 28051 sw
rect 30064 28035 30173 28043
tri 30173 28035 30181 28043 sw
rect 30064 28027 30181 28035
tri 30181 28027 30189 28035 sw
rect 30064 28019 30189 28027
tri 30189 28019 30197 28027 sw
rect 30064 28014 30197 28019
rect 29929 28011 30197 28014
tri 30197 28011 30205 28019 sw
tri 29929 28003 29937 28011 ne
rect 29937 28003 30205 28011
tri 30205 28003 30213 28011 sw
tri 29937 27995 29945 28003 ne
rect 29945 27995 30213 28003
tri 30213 27995 30221 28003 sw
rect 70802 27996 71000 28054
tri 29945 27992 29948 27995 ne
rect 29948 27992 30221 27995
tri 29948 27984 29956 27992 ne
rect 29956 27987 30221 27992
tri 30221 27987 30229 27995 sw
rect 29956 27984 30229 27987
tri 29956 27976 29964 27984 ne
rect 29964 27979 30229 27984
tri 30229 27979 30237 27987 sw
rect 29964 27976 30237 27979
tri 29964 27968 29972 27976 ne
rect 29972 27971 30237 27976
tri 30237 27971 30245 27979 sw
rect 29972 27968 30245 27971
tri 29972 27960 29980 27968 ne
rect 29980 27963 30245 27968
tri 30245 27963 30253 27971 sw
rect 29980 27960 30253 27963
tri 29980 27952 29988 27960 ne
rect 29988 27955 30253 27960
tri 30253 27955 30261 27963 sw
rect 29988 27952 30261 27955
tri 29988 27944 29996 27952 ne
rect 29996 27947 30261 27952
tri 30261 27947 30269 27955 sw
rect 70802 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 29996 27944 30269 27947
tri 29996 27936 30004 27944 ne
rect 30004 27939 30269 27944
tri 30269 27939 30277 27947 sw
rect 30004 27936 30277 27939
tri 30004 27928 30012 27936 ne
rect 30012 27931 30277 27936
tri 30277 27931 30285 27939 sw
rect 30012 27928 30285 27931
tri 30012 27920 30020 27928 ne
rect 30020 27920 30150 27928
tri 30020 27912 30028 27920 ne
rect 30028 27912 30150 27920
tri 30028 27904 30036 27912 ne
rect 30036 27904 30150 27912
tri 30036 27896 30044 27904 ne
rect 30044 27896 30150 27904
tri 30044 27888 30052 27896 ne
rect 30052 27888 30150 27896
tri 30052 27880 30060 27888 ne
rect 30060 27882 30150 27888
rect 30196 27923 30285 27928
tri 30285 27923 30293 27931 sw
rect 30196 27919 30293 27923
tri 30293 27919 30297 27923 sw
rect 30196 27911 30297 27919
tri 30297 27911 30305 27919 sw
rect 30196 27903 30305 27911
tri 30305 27903 30313 27911 sw
rect 30196 27895 30313 27903
tri 30313 27895 30321 27903 sw
rect 30196 27887 30321 27895
tri 30321 27887 30329 27895 sw
rect 70802 27892 71000 27950
rect 30196 27882 30329 27887
rect 30060 27880 30329 27882
tri 30060 27879 30061 27880 ne
rect 30061 27879 30329 27880
tri 30329 27879 30337 27887 sw
tri 30061 27871 30069 27879 ne
rect 30069 27871 30337 27879
tri 30337 27871 30345 27879 sw
tri 30069 27863 30077 27871 ne
rect 30077 27863 30345 27871
tri 30345 27863 30353 27871 sw
tri 30077 27855 30085 27863 ne
rect 30085 27855 30353 27863
tri 30353 27855 30361 27863 sw
tri 30085 27847 30093 27855 ne
rect 30093 27847 30361 27855
tri 30361 27847 30369 27855 sw
tri 30093 27839 30101 27847 ne
rect 30101 27839 30369 27847
tri 30369 27839 30377 27847 sw
rect 70802 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30101 27831 30109 27839 ne
rect 30109 27831 30377 27839
tri 30377 27831 30385 27839 sw
tri 30109 27823 30117 27831 ne
rect 30117 27823 30385 27831
tri 30385 27823 30393 27831 sw
tri 30117 27815 30125 27823 ne
rect 30125 27815 30393 27823
tri 30393 27815 30401 27823 sw
tri 30125 27807 30133 27815 ne
rect 30133 27807 30401 27815
tri 30401 27807 30409 27815 sw
tri 30133 27799 30141 27807 ne
rect 30141 27799 30409 27807
tri 30409 27799 30417 27807 sw
tri 30141 27795 30145 27799 ne
rect 30145 27796 30417 27799
rect 30145 27795 30282 27796
tri 30145 27791 30149 27795 ne
rect 30149 27791 30282 27795
tri 30149 27783 30157 27791 ne
rect 30157 27783 30282 27791
tri 30157 27775 30165 27783 ne
rect 30165 27775 30282 27783
tri 30165 27767 30173 27775 ne
rect 30173 27767 30282 27775
tri 30173 27759 30181 27767 ne
rect 30181 27759 30282 27767
tri 30181 27751 30189 27759 ne
rect 30189 27751 30282 27759
tri 30189 27743 30197 27751 ne
rect 30197 27750 30282 27751
rect 30328 27791 30417 27796
tri 30417 27791 30425 27799 sw
rect 30328 27783 30425 27791
tri 30425 27783 30433 27791 sw
rect 70802 27788 71000 27846
rect 30328 27775 30433 27783
tri 30433 27775 30441 27783 sw
rect 30328 27767 30441 27775
tri 30441 27767 30449 27775 sw
rect 30328 27759 30449 27767
tri 30449 27759 30457 27767 sw
rect 30328 27751 30457 27759
tri 30457 27751 30465 27759 sw
rect 30328 27750 30465 27751
rect 30197 27745 30465 27750
tri 30465 27745 30471 27751 sw
rect 30197 27743 30471 27745
tri 30197 27735 30205 27743 ne
rect 30205 27737 30471 27743
tri 30471 27737 30479 27745 sw
rect 70802 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
rect 30205 27735 30479 27737
tri 30205 27727 30213 27735 ne
rect 30213 27729 30479 27735
tri 30479 27729 30487 27737 sw
rect 30213 27727 30487 27729
tri 30213 27724 30216 27727 ne
rect 30216 27724 30487 27727
tri 30216 27716 30224 27724 ne
rect 30224 27721 30487 27724
tri 30487 27721 30495 27729 sw
rect 30224 27716 30495 27721
tri 30224 27708 30232 27716 ne
rect 30232 27713 30495 27716
tri 30495 27713 30503 27721 sw
rect 30232 27708 30503 27713
tri 30232 27700 30240 27708 ne
rect 30240 27705 30503 27708
tri 30503 27705 30511 27713 sw
rect 30240 27700 30511 27705
tri 30240 27692 30248 27700 ne
rect 30248 27697 30511 27700
tri 30511 27697 30519 27705 sw
rect 30248 27692 30519 27697
tri 30248 27684 30256 27692 ne
rect 30256 27689 30519 27692
tri 30519 27689 30527 27697 sw
rect 30256 27684 30527 27689
tri 30256 27676 30264 27684 ne
rect 30264 27681 30527 27684
tri 30527 27681 30535 27689 sw
rect 70802 27684 71000 27742
rect 30264 27676 30535 27681
tri 30264 27668 30272 27676 ne
rect 30272 27673 30535 27676
tri 30535 27673 30543 27681 sw
rect 30272 27668 30543 27673
tri 30272 27660 30280 27668 ne
rect 30280 27665 30543 27668
tri 30543 27665 30551 27673 sw
rect 30280 27664 30551 27665
rect 30280 27660 30414 27664
tri 30280 27652 30288 27660 ne
rect 30288 27652 30414 27660
tri 30288 27644 30296 27652 ne
rect 30296 27644 30414 27652
tri 30296 27636 30304 27644 ne
rect 30304 27636 30414 27644
tri 30304 27628 30312 27636 ne
rect 30312 27628 30414 27636
tri 30312 27620 30320 27628 ne
rect 30320 27620 30414 27628
tri 30320 27612 30328 27620 ne
rect 30328 27618 30414 27620
rect 30460 27657 30551 27664
tri 30551 27657 30559 27665 sw
rect 30460 27649 30559 27657
tri 30559 27649 30567 27657 sw
rect 30460 27641 30567 27649
tri 30567 27641 30575 27649 sw
rect 30460 27633 30575 27641
tri 30575 27633 30583 27641 sw
rect 70802 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30460 27625 30583 27633
tri 30583 27625 30591 27633 sw
rect 30460 27619 30591 27625
tri 30591 27619 30597 27625 sw
rect 30460 27618 30597 27619
rect 30328 27612 30597 27618
tri 30328 27604 30336 27612 ne
rect 30336 27611 30597 27612
tri 30597 27611 30605 27619 sw
rect 30336 27604 30605 27611
tri 30336 27596 30344 27604 ne
rect 30344 27603 30605 27604
tri 30605 27603 30613 27611 sw
rect 30344 27596 30613 27603
tri 30344 27590 30350 27596 ne
rect 30350 27595 30613 27596
tri 30613 27595 30621 27603 sw
rect 30350 27590 30621 27595
tri 30350 27582 30358 27590 ne
rect 30358 27587 30621 27590
tri 30621 27587 30629 27595 sw
rect 30358 27582 30629 27587
tri 30358 27574 30366 27582 ne
rect 30366 27579 30629 27582
tri 30629 27579 30637 27587 sw
rect 70802 27580 71000 27638
rect 30366 27574 30637 27579
tri 30366 27566 30374 27574 ne
rect 30374 27571 30637 27574
tri 30637 27571 30645 27579 sw
rect 30374 27566 30645 27571
tri 30374 27558 30382 27566 ne
rect 30382 27563 30645 27566
tri 30645 27563 30653 27571 sw
rect 30382 27558 30653 27563
tri 30382 27550 30390 27558 ne
rect 30390 27555 30653 27558
tri 30653 27555 30661 27563 sw
rect 30390 27550 30661 27555
tri 30390 27542 30398 27550 ne
rect 30398 27547 30661 27550
tri 30661 27547 30669 27555 sw
rect 30398 27542 30669 27547
tri 30398 27534 30406 27542 ne
rect 30406 27539 30669 27542
tri 30669 27539 30677 27547 sw
rect 30406 27534 30677 27539
tri 30406 27526 30414 27534 ne
rect 30414 27532 30677 27534
rect 30414 27526 30546 27532
tri 30414 27523 30417 27526 ne
rect 30417 27523 30546 27526
tri 30417 27515 30425 27523 ne
rect 30425 27515 30546 27523
tri 30425 27507 30433 27515 ne
rect 30433 27507 30546 27515
tri 30433 27499 30441 27507 ne
rect 30441 27499 30546 27507
tri 30441 27491 30449 27499 ne
rect 30449 27491 30546 27499
tri 30449 27483 30457 27491 ne
rect 30457 27486 30546 27491
rect 30592 27531 30677 27532
tri 30677 27531 30685 27539 sw
rect 70802 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 30592 27523 30685 27531
tri 30685 27523 30693 27531 sw
rect 30592 27515 30693 27523
tri 30693 27515 30701 27523 sw
rect 30592 27507 30701 27515
tri 30701 27507 30709 27515 sw
rect 30592 27499 30709 27507
tri 30709 27499 30717 27507 sw
rect 30592 27491 30717 27499
tri 30717 27491 30725 27499 sw
rect 30592 27486 30725 27491
rect 30457 27483 30725 27486
tri 30725 27483 30733 27491 sw
tri 30457 27475 30465 27483 ne
rect 30465 27475 30733 27483
tri 30733 27475 30741 27483 sw
rect 70802 27476 71000 27534
tri 30465 27467 30473 27475 ne
rect 30473 27467 30741 27475
tri 30741 27467 30749 27475 sw
tri 30473 27459 30481 27467 ne
rect 30481 27459 30749 27467
tri 30749 27459 30757 27467 sw
tri 30481 27452 30488 27459 ne
rect 30488 27452 30757 27459
tri 30757 27452 30764 27459 sw
tri 30488 27444 30496 27452 ne
rect 30496 27444 30764 27452
tri 30764 27444 30772 27452 sw
tri 30496 27436 30504 27444 ne
rect 30504 27436 30772 27444
tri 30772 27436 30780 27444 sw
tri 30504 27428 30512 27436 ne
rect 30512 27428 30780 27436
tri 30780 27428 30788 27436 sw
rect 70802 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30512 27420 30520 27428 ne
rect 30520 27420 30788 27428
tri 30788 27420 30796 27428 sw
tri 30520 27412 30528 27420 ne
rect 30528 27412 30796 27420
tri 30796 27412 30804 27420 sw
tri 30528 27404 30536 27412 ne
rect 30536 27404 30804 27412
tri 30804 27404 30812 27412 sw
tri 30536 27396 30544 27404 ne
rect 30544 27400 30812 27404
rect 30544 27396 30678 27400
tri 30544 27388 30552 27396 ne
rect 30552 27388 30678 27396
tri 30552 27380 30560 27388 ne
rect 30560 27380 30678 27388
tri 30560 27372 30568 27380 ne
rect 30568 27372 30678 27380
tri 30568 27364 30576 27372 ne
rect 30576 27364 30678 27372
tri 30576 27356 30584 27364 ne
rect 30584 27356 30678 27364
tri 30584 27348 30592 27356 ne
rect 30592 27354 30678 27356
rect 30724 27396 30812 27400
tri 30812 27396 30820 27404 sw
rect 30724 27388 30820 27396
tri 30820 27388 30828 27396 sw
rect 30724 27380 30828 27388
tri 30828 27380 30836 27388 sw
rect 30724 27372 30836 27380
tri 30836 27372 30844 27380 sw
rect 70802 27372 71000 27430
rect 30724 27364 30844 27372
tri 30844 27364 30852 27372 sw
rect 30724 27356 30852 27364
tri 30852 27356 30860 27364 sw
rect 30724 27354 30860 27356
rect 30592 27348 30860 27354
tri 30860 27348 30868 27356 sw
tri 30592 27340 30600 27348 ne
rect 30600 27343 30868 27348
tri 30868 27343 30873 27348 sw
rect 30600 27340 30873 27343
tri 30600 27332 30608 27340 ne
rect 30608 27335 30873 27340
tri 30873 27335 30881 27343 sw
rect 30608 27332 30881 27335
tri 30608 27330 30610 27332 ne
rect 30610 27330 30881 27332
tri 30610 27322 30618 27330 ne
rect 30618 27327 30881 27330
tri 30881 27327 30889 27335 sw
rect 30618 27322 30889 27327
tri 30618 27314 30626 27322 ne
rect 30626 27319 30889 27322
tri 30889 27319 30897 27327 sw
rect 70802 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
rect 30626 27314 30897 27319
tri 30626 27306 30634 27314 ne
rect 30634 27311 30897 27314
tri 30897 27311 30905 27319 sw
rect 30634 27306 30905 27311
tri 30634 27298 30642 27306 ne
rect 30642 27303 30905 27306
tri 30905 27303 30913 27311 sw
rect 30642 27298 30913 27303
tri 30642 27290 30650 27298 ne
rect 30650 27295 30913 27298
tri 30913 27295 30921 27303 sw
rect 30650 27290 30921 27295
tri 30650 27282 30658 27290 ne
rect 30658 27287 30921 27290
tri 30921 27287 30929 27295 sw
rect 30658 27282 30929 27287
tri 30658 27274 30666 27282 ne
rect 30666 27279 30929 27282
tri 30929 27279 30937 27287 sw
rect 30666 27274 30937 27279
tri 30666 27266 30674 27274 ne
rect 30674 27271 30937 27274
tri 30937 27271 30945 27279 sw
rect 30674 27268 30945 27271
rect 30674 27266 30810 27268
tri 30674 27258 30682 27266 ne
rect 30682 27258 30810 27266
tri 30682 27250 30690 27258 ne
rect 30690 27250 30810 27258
tri 30690 27242 30698 27250 ne
rect 30698 27242 30810 27250
tri 30698 27234 30706 27242 ne
rect 30706 27234 30810 27242
tri 30706 27226 30714 27234 ne
rect 30714 27226 30810 27234
tri 30714 27218 30722 27226 ne
rect 30722 27222 30810 27226
rect 30856 27266 30945 27268
tri 30945 27266 30950 27271 sw
rect 70802 27268 71000 27326
rect 30856 27258 30950 27266
tri 30950 27258 30958 27266 sw
rect 30856 27250 30958 27258
tri 30958 27250 30966 27258 sw
rect 30856 27242 30966 27250
tri 30966 27242 30974 27250 sw
rect 30856 27234 30974 27242
tri 30974 27234 30982 27242 sw
rect 30856 27226 30982 27234
tri 30982 27226 30990 27234 sw
rect 30856 27222 30990 27226
rect 30722 27218 30990 27222
tri 30990 27218 30998 27226 sw
rect 70802 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30722 27213 30727 27218 ne
rect 30727 27213 30998 27218
tri 30998 27213 31003 27218 sw
tri 30727 27205 30735 27213 ne
rect 30735 27205 31003 27213
tri 31003 27205 31011 27213 sw
tri 30735 27197 30743 27205 ne
rect 30743 27197 31011 27205
tri 31011 27197 31019 27205 sw
tri 30743 27189 30751 27197 ne
rect 30751 27189 31019 27197
tri 31019 27189 31027 27197 sw
tri 30751 27181 30759 27189 ne
rect 30759 27181 31027 27189
tri 31027 27181 31035 27189 sw
tri 30759 27173 30767 27181 ne
rect 30767 27173 31035 27181
tri 31035 27173 31043 27181 sw
tri 30767 27165 30775 27173 ne
rect 30775 27165 31043 27173
tri 31043 27165 31051 27173 sw
tri 30775 27157 30783 27165 ne
rect 30783 27157 31051 27165
tri 31051 27157 31059 27165 sw
rect 70802 27164 71000 27222
tri 30783 27149 30791 27157 ne
rect 30791 27149 31059 27157
tri 31059 27149 31067 27157 sw
tri 30791 27141 30799 27149 ne
rect 30799 27141 31067 27149
tri 31067 27141 31075 27149 sw
tri 30799 27133 30807 27141 ne
rect 30807 27136 31075 27141
rect 30807 27133 30942 27136
tri 30807 27125 30815 27133 ne
rect 30815 27125 30942 27133
tri 30815 27117 30823 27125 ne
rect 30823 27117 30942 27125
tri 30823 27109 30831 27117 ne
rect 30831 27109 30942 27117
tri 30831 27101 30839 27109 ne
rect 30839 27101 30942 27109
tri 30839 27093 30847 27101 ne
rect 30847 27093 30942 27101
tri 30847 27085 30855 27093 ne
rect 30855 27090 30942 27093
rect 30988 27133 31075 27136
tri 31075 27133 31083 27141 sw
rect 30988 27125 31083 27133
tri 31083 27125 31091 27133 sw
rect 30988 27117 31091 27125
tri 31091 27117 31099 27125 sw
rect 70802 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 30988 27109 31099 27117
tri 31099 27109 31107 27117 sw
rect 30988 27101 31107 27109
tri 31107 27101 31115 27109 sw
rect 30988 27098 31115 27101
tri 31115 27098 31118 27101 sw
rect 30988 27090 31118 27098
tri 31118 27090 31126 27098 sw
rect 30855 27085 31126 27090
tri 30855 27083 30857 27085 ne
rect 30857 27083 31126 27085
tri 30857 27075 30865 27083 ne
rect 30865 27082 31126 27083
tri 31126 27082 31134 27090 sw
rect 30865 27075 31134 27082
tri 30865 27067 30873 27075 ne
rect 30873 27074 31134 27075
tri 31134 27074 31142 27082 sw
rect 30873 27067 31142 27074
tri 30873 27059 30881 27067 ne
rect 30881 27066 31142 27067
tri 31142 27066 31150 27074 sw
rect 30881 27059 31150 27066
tri 30881 27051 30889 27059 ne
rect 30889 27058 31150 27059
tri 31150 27058 31158 27066 sw
rect 70802 27060 71000 27118
rect 30889 27051 31158 27058
tri 30889 27043 30897 27051 ne
rect 30897 27050 31158 27051
tri 31158 27050 31166 27058 sw
rect 30897 27043 31166 27050
tri 30897 27035 30905 27043 ne
rect 30905 27042 31166 27043
tri 31166 27042 31174 27050 sw
rect 30905 27035 31174 27042
tri 30905 27027 30913 27035 ne
rect 30913 27034 31174 27035
tri 31174 27034 31182 27042 sw
rect 30913 27027 31182 27034
tri 30913 27019 30921 27027 ne
rect 30921 27026 31182 27027
tri 31182 27026 31190 27034 sw
rect 30921 27019 31190 27026
tri 30921 27011 30929 27019 ne
rect 30929 27018 31190 27019
tri 31190 27018 31198 27026 sw
rect 30929 27011 31198 27018
tri 30929 27003 30937 27011 ne
rect 30937 27010 31198 27011
tri 31198 27010 31206 27018 sw
rect 70802 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 30937 27004 31206 27010
rect 30937 27003 31074 27004
tri 30937 26998 30942 27003 ne
rect 30942 26998 31074 27003
tri 30942 26995 30945 26998 ne
rect 30945 26995 31074 26998
tri 30945 26987 30953 26995 ne
rect 30953 26987 31074 26995
tri 30953 26979 30961 26987 ne
rect 30961 26979 31074 26987
tri 30961 26971 30969 26979 ne
rect 30969 26971 31074 26979
tri 30969 26963 30977 26971 ne
rect 30977 26963 31074 26971
tri 30977 26955 30985 26963 ne
rect 30985 26958 31074 26963
rect 31120 27003 31206 27004
tri 31206 27003 31213 27010 sw
rect 31120 26995 31213 27003
tri 31213 26995 31221 27003 sw
rect 31120 26987 31221 26995
tri 31221 26987 31229 26995 sw
rect 31120 26979 31229 26987
tri 31229 26979 31237 26987 sw
rect 31120 26971 31237 26979
tri 31237 26971 31245 26979 sw
rect 31120 26963 31245 26971
tri 31245 26963 31253 26971 sw
rect 31120 26958 31253 26963
rect 30985 26955 31253 26958
tri 31253 26955 31261 26963 sw
rect 70802 26956 71000 27014
tri 30985 26947 30993 26955 ne
rect 30993 26947 31261 26955
tri 31261 26947 31269 26955 sw
tri 30993 26939 31001 26947 ne
rect 31001 26945 31269 26947
tri 31269 26945 31271 26947 sw
rect 31001 26939 31271 26945
tri 31001 26931 31009 26939 ne
rect 31009 26937 31271 26939
tri 31271 26937 31279 26945 sw
rect 31009 26931 31279 26937
tri 31009 26930 31010 26931 ne
rect 31010 26930 31279 26931
tri 31010 26922 31018 26930 ne
rect 31018 26929 31279 26930
tri 31279 26929 31287 26937 sw
rect 31018 26922 31287 26929
tri 31018 26914 31026 26922 ne
rect 31026 26921 31287 26922
tri 31287 26921 31295 26929 sw
rect 31026 26914 31295 26921
tri 31026 26906 31034 26914 ne
rect 31034 26913 31295 26914
tri 31295 26913 31303 26921 sw
rect 31034 26906 31303 26913
tri 31034 26898 31042 26906 ne
rect 31042 26905 31303 26906
tri 31303 26905 31311 26913 sw
rect 70802 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
rect 31042 26898 31311 26905
tri 31042 26890 31050 26898 ne
rect 31050 26897 31311 26898
tri 31311 26897 31319 26905 sw
rect 31050 26890 31319 26897
tri 31050 26882 31058 26890 ne
rect 31058 26889 31319 26890
tri 31319 26889 31327 26897 sw
rect 31058 26882 31327 26889
tri 31058 26874 31066 26882 ne
rect 31066 26881 31327 26882
tri 31327 26881 31335 26889 sw
rect 31066 26874 31335 26881
tri 31066 26866 31074 26874 ne
rect 31074 26873 31335 26874
tri 31335 26873 31343 26881 sw
rect 31074 26872 31343 26873
rect 31074 26866 31206 26872
tri 31074 26858 31082 26866 ne
rect 31082 26858 31206 26866
tri 31082 26850 31090 26858 ne
rect 31090 26850 31206 26858
tri 31090 26842 31098 26850 ne
rect 31098 26842 31206 26850
tri 31098 26834 31106 26842 ne
rect 31106 26834 31206 26842
tri 31106 26826 31114 26834 ne
rect 31114 26826 31206 26834
rect 31252 26865 31343 26872
tri 31343 26865 31351 26873 sw
rect 31252 26857 31351 26865
tri 31351 26857 31359 26865 sw
rect 31252 26849 31359 26857
tri 31359 26849 31367 26857 sw
rect 70802 26852 71000 26910
rect 31252 26841 31367 26849
tri 31367 26841 31375 26849 sw
rect 31252 26833 31375 26841
tri 31375 26833 31383 26841 sw
rect 31252 26832 31383 26833
tri 31383 26832 31384 26833 sw
rect 31252 26826 31384 26832
tri 31114 26818 31122 26826 ne
rect 31122 26824 31384 26826
tri 31384 26824 31392 26832 sw
rect 31122 26818 31392 26824
tri 31122 26810 31130 26818 ne
rect 31130 26816 31392 26818
tri 31392 26816 31400 26824 sw
rect 31130 26810 31400 26816
tri 31130 26802 31138 26810 ne
rect 31138 26808 31400 26810
tri 31400 26808 31408 26816 sw
rect 31138 26802 31408 26808
tri 31138 26794 31146 26802 ne
rect 31146 26800 31408 26802
tri 31408 26800 31416 26808 sw
rect 70802 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 31146 26794 31416 26800
tri 31146 26786 31154 26794 ne
rect 31154 26792 31416 26794
tri 31416 26792 31424 26800 sw
rect 31154 26786 31424 26792
tri 31154 26778 31162 26786 ne
rect 31162 26784 31424 26786
tri 31424 26784 31432 26792 sw
rect 31162 26778 31432 26784
tri 31162 26770 31170 26778 ne
rect 31170 26776 31432 26778
tri 31432 26776 31440 26784 sw
rect 31170 26770 31440 26776
tri 31170 26762 31178 26770 ne
rect 31178 26768 31440 26770
tri 31440 26768 31448 26776 sw
rect 31178 26762 31448 26768
tri 31178 26754 31186 26762 ne
rect 31186 26760 31448 26762
tri 31448 26760 31456 26768 sw
rect 31186 26756 31456 26760
tri 31456 26756 31460 26760 sw
rect 31186 26754 31460 26756
tri 31186 26746 31194 26754 ne
rect 31194 26752 31460 26754
tri 31460 26752 31464 26756 sw
rect 31194 26746 31464 26752
tri 31194 26738 31202 26746 ne
rect 31202 26744 31464 26746
tri 31464 26744 31472 26752 sw
rect 70802 26748 71000 26806
rect 31202 26740 31472 26744
rect 31202 26738 31338 26740
tri 31202 26734 31206 26738 ne
rect 31206 26734 31338 26738
tri 31206 26730 31210 26734 ne
rect 31210 26730 31338 26734
tri 31210 26722 31218 26730 ne
rect 31218 26722 31338 26730
tri 31218 26714 31226 26722 ne
rect 31226 26714 31338 26722
tri 31226 26706 31234 26714 ne
rect 31234 26706 31338 26714
tri 31234 26698 31242 26706 ne
rect 31242 26698 31338 26706
tri 31242 26690 31250 26698 ne
rect 31250 26694 31338 26698
rect 31384 26736 31472 26740
tri 31472 26736 31480 26744 sw
rect 31384 26728 31480 26736
tri 31480 26728 31488 26736 sw
rect 31384 26720 31488 26728
tri 31488 26720 31496 26728 sw
rect 31384 26712 31496 26720
tri 31496 26712 31504 26720 sw
rect 31384 26704 31504 26712
tri 31504 26704 31512 26712 sw
rect 31384 26696 31512 26704
tri 31512 26696 31520 26704 sw
rect 70802 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 31384 26694 31520 26696
rect 31250 26690 31520 26694
tri 31250 26682 31258 26690 ne
rect 31258 26688 31520 26690
tri 31520 26688 31528 26696 sw
rect 31258 26682 31528 26688
tri 31258 26674 31266 26682 ne
rect 31266 26680 31528 26682
tri 31528 26680 31536 26688 sw
rect 31266 26674 31536 26680
tri 31266 26666 31274 26674 ne
rect 31274 26672 31536 26674
tri 31536 26672 31544 26680 sw
rect 31274 26666 31544 26672
tri 31274 26658 31282 26666 ne
rect 31282 26664 31544 26666
tri 31544 26664 31552 26672 sw
rect 31282 26658 31552 26664
tri 31282 26650 31290 26658 ne
rect 31290 26656 31552 26658
tri 31552 26656 31560 26664 sw
rect 31290 26650 31560 26656
tri 31290 26642 31298 26650 ne
rect 31298 26648 31560 26650
tri 31560 26648 31568 26656 sw
rect 31298 26642 31568 26648
tri 31298 26634 31306 26642 ne
rect 31306 26640 31568 26642
tri 31568 26640 31576 26648 sw
rect 70802 26644 71000 26702
rect 31306 26637 31576 26640
tri 31576 26637 31579 26640 sw
rect 31306 26634 31579 26637
tri 31306 26626 31314 26634 ne
rect 31314 26629 31579 26634
tri 31579 26629 31587 26637 sw
rect 31314 26626 31587 26629
tri 31314 26618 31322 26626 ne
rect 31322 26621 31587 26626
tri 31587 26621 31595 26629 sw
rect 31322 26618 31595 26621
tri 31322 26613 31327 26618 ne
rect 31327 26613 31595 26618
tri 31595 26613 31603 26621 sw
tri 31327 26605 31335 26613 ne
rect 31335 26608 31603 26613
rect 31335 26605 31470 26608
tri 31335 26597 31343 26605 ne
rect 31343 26597 31470 26605
tri 31343 26589 31351 26597 ne
rect 31351 26589 31470 26597
tri 31351 26581 31359 26589 ne
rect 31359 26581 31470 26589
tri 31359 26573 31367 26581 ne
rect 31367 26573 31470 26581
tri 31367 26565 31375 26573 ne
rect 31375 26565 31470 26573
tri 31375 26557 31383 26565 ne
rect 31383 26562 31470 26565
rect 31516 26605 31603 26608
tri 31603 26605 31611 26613 sw
rect 31516 26597 31611 26605
tri 31611 26597 31619 26605 sw
rect 70802 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 31516 26589 31619 26597
tri 31619 26589 31627 26597 sw
rect 31516 26581 31627 26589
tri 31627 26581 31635 26589 sw
rect 31516 26573 31635 26581
tri 31635 26573 31643 26581 sw
rect 31516 26565 31643 26573
tri 31643 26565 31651 26573 sw
rect 31516 26562 31651 26565
rect 31383 26557 31651 26562
tri 31651 26557 31659 26565 sw
tri 31383 26549 31391 26557 ne
rect 31391 26549 31659 26557
tri 31659 26549 31667 26557 sw
tri 31391 26541 31399 26549 ne
rect 31399 26541 31667 26549
tri 31667 26541 31675 26549 sw
tri 31399 26533 31407 26541 ne
rect 31407 26533 31675 26541
tri 31675 26533 31683 26541 sw
rect 70802 26540 71000 26598
tri 31407 26525 31415 26533 ne
rect 31415 26525 31683 26533
tri 31683 26525 31691 26533 sw
tri 31415 26517 31423 26525 ne
rect 31423 26517 31691 26525
tri 31691 26517 31699 26525 sw
tri 31423 26509 31431 26517 ne
rect 31431 26509 31699 26517
tri 31699 26509 31707 26517 sw
tri 31431 26501 31439 26509 ne
rect 31439 26501 31707 26509
tri 31707 26501 31715 26509 sw
tri 31439 26493 31447 26501 ne
rect 31447 26499 31715 26501
tri 31715 26499 31717 26501 sw
rect 31447 26493 31717 26499
tri 31447 26491 31449 26493 ne
rect 31449 26491 31717 26493
tri 31717 26491 31725 26499 sw
rect 70802 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
tri 31449 26483 31457 26491 ne
rect 31457 26483 31725 26491
tri 31725 26483 31733 26491 sw
tri 31457 26476 31464 26483 ne
rect 31464 26476 31733 26483
tri 31464 26475 31465 26476 ne
rect 31465 26475 31602 26476
tri 31465 26467 31473 26475 ne
rect 31473 26467 31602 26475
tri 31473 26459 31481 26467 ne
rect 31481 26459 31602 26467
tri 31481 26451 31489 26459 ne
rect 31489 26451 31602 26459
tri 31489 26443 31497 26451 ne
rect 31497 26443 31602 26451
tri 31497 26435 31505 26443 ne
rect 31505 26435 31602 26443
tri 31505 26427 31513 26435 ne
rect 31513 26430 31602 26435
rect 31648 26475 31733 26476
tri 31733 26475 31741 26483 sw
rect 31648 26467 31741 26475
tri 31741 26467 31749 26475 sw
rect 31648 26459 31749 26467
tri 31749 26459 31757 26467 sw
rect 31648 26451 31757 26459
tri 31757 26451 31765 26459 sw
rect 31648 26443 31765 26451
tri 31765 26443 31773 26451 sw
rect 31648 26435 31773 26443
tri 31773 26435 31781 26443 sw
rect 70802 26436 71000 26494
rect 31648 26430 31781 26435
rect 31513 26427 31781 26430
tri 31781 26427 31789 26435 sw
tri 31513 26419 31521 26427 ne
rect 31521 26419 31789 26427
tri 31789 26419 31797 26427 sw
tri 31521 26411 31529 26419 ne
rect 31529 26411 31797 26419
tri 31797 26411 31805 26419 sw
tri 31529 26403 31537 26411 ne
rect 31537 26403 31805 26411
tri 31805 26403 31813 26411 sw
tri 31537 26395 31545 26403 ne
rect 31545 26395 31813 26403
tri 31813 26395 31821 26403 sw
tri 31545 26387 31553 26395 ne
rect 31553 26387 31821 26395
tri 31821 26387 31829 26395 sw
rect 70802 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31553 26379 31561 26387 ne
rect 31561 26379 31829 26387
tri 31829 26379 31837 26387 sw
tri 31561 26371 31569 26379 ne
rect 31569 26371 31837 26379
tri 31837 26371 31845 26379 sw
tri 31569 26363 31577 26371 ne
rect 31577 26363 31845 26371
tri 31845 26363 31853 26371 sw
tri 31577 26355 31585 26363 ne
rect 31585 26357 31853 26363
tri 31853 26357 31859 26363 sw
rect 31585 26355 31859 26357
tri 31585 26353 31587 26355 ne
rect 31587 26353 31859 26355
tri 31587 26345 31595 26353 ne
rect 31595 26349 31859 26353
tri 31859 26349 31867 26357 sw
rect 31595 26345 31867 26349
tri 31595 26337 31603 26345 ne
rect 31603 26344 31867 26345
rect 31603 26337 31734 26344
tri 31603 26329 31611 26337 ne
rect 31611 26329 31734 26337
tri 31611 26321 31619 26329 ne
rect 31619 26321 31734 26329
tri 31619 26313 31627 26321 ne
rect 31627 26313 31734 26321
tri 31627 26305 31635 26313 ne
rect 31635 26305 31734 26313
tri 31635 26297 31643 26305 ne
rect 31643 26298 31734 26305
rect 31780 26341 31867 26344
tri 31867 26341 31875 26349 sw
rect 31780 26333 31875 26341
tri 31875 26333 31883 26341 sw
rect 31780 26325 31883 26333
tri 31883 26325 31891 26333 sw
rect 70802 26332 71000 26390
rect 31780 26317 31891 26325
tri 31891 26317 31899 26325 sw
rect 31780 26309 31899 26317
tri 31899 26309 31907 26317 sw
rect 31780 26301 31907 26309
tri 31907 26301 31915 26309 sw
rect 31780 26298 31915 26301
rect 31643 26297 31915 26298
tri 31643 26289 31651 26297 ne
rect 31651 26293 31915 26297
tri 31915 26293 31923 26301 sw
rect 31651 26289 31923 26293
tri 31651 26281 31659 26289 ne
rect 31659 26285 31923 26289
tri 31923 26285 31931 26293 sw
rect 70802 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
rect 31659 26281 31931 26285
tri 31659 26273 31667 26281 ne
rect 31667 26277 31931 26281
tri 31931 26277 31939 26285 sw
rect 31667 26273 31939 26277
tri 31667 26265 31675 26273 ne
rect 31675 26269 31939 26273
tri 31939 26269 31947 26277 sw
rect 31675 26265 31947 26269
tri 31675 26257 31683 26265 ne
rect 31683 26261 31947 26265
tri 31947 26261 31955 26269 sw
rect 31683 26257 31955 26261
tri 31683 26249 31691 26257 ne
rect 31691 26253 31955 26257
tri 31955 26253 31963 26261 sw
rect 31691 26249 31963 26253
tri 31691 26241 31699 26249 ne
rect 31699 26245 31963 26249
tri 31963 26245 31971 26253 sw
rect 31699 26241 31971 26245
tri 31971 26241 31975 26245 sw
tri 31699 26239 31701 26241 ne
rect 31701 26239 31975 26241
tri 31701 26231 31709 26239 ne
rect 31709 26237 31975 26239
tri 31975 26237 31979 26241 sw
rect 31709 26231 31979 26237
tri 31979 26231 31985 26237 sw
tri 31709 26223 31717 26231 ne
rect 31717 26223 31985 26231
tri 31985 26223 31993 26231 sw
rect 70802 26228 71000 26286
tri 31717 26215 31725 26223 ne
rect 31725 26215 31993 26223
tri 31993 26215 32001 26223 sw
tri 31725 26207 31733 26215 ne
rect 31733 26212 32001 26215
rect 31733 26207 31866 26212
tri 31733 26199 31741 26207 ne
rect 31741 26199 31866 26207
tri 31741 26191 31749 26199 ne
rect 31749 26191 31866 26199
tri 31749 26183 31757 26191 ne
rect 31757 26183 31866 26191
tri 31757 26175 31765 26183 ne
rect 31765 26175 31866 26183
tri 31765 26167 31773 26175 ne
rect 31773 26167 31866 26175
tri 31773 26159 31781 26167 ne
rect 31781 26166 31866 26167
rect 31912 26207 32001 26212
tri 32001 26207 32009 26215 sw
rect 31912 26199 32009 26207
tri 32009 26199 32017 26207 sw
rect 31912 26191 32017 26199
tri 32017 26191 32025 26199 sw
rect 31912 26183 32025 26191
tri 32025 26183 32033 26191 sw
rect 31912 26175 32033 26183
tri 32033 26175 32041 26183 sw
rect 70802 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 31912 26170 32041 26175
tri 32041 26170 32046 26175 sw
rect 31912 26166 32046 26170
rect 31781 26162 32046 26166
tri 32046 26162 32054 26170 sw
rect 31781 26159 32054 26162
tri 31781 26151 31789 26159 ne
rect 31789 26154 32054 26159
tri 32054 26154 32062 26162 sw
rect 31789 26151 32062 26154
tri 31789 26143 31797 26151 ne
rect 31797 26146 32062 26151
tri 32062 26146 32070 26154 sw
rect 31797 26143 32070 26146
tri 31797 26135 31805 26143 ne
rect 31805 26138 32070 26143
tri 32070 26138 32078 26146 sw
rect 31805 26135 32078 26138
tri 31805 26127 31813 26135 ne
rect 31813 26130 32078 26135
tri 32078 26130 32086 26138 sw
rect 31813 26127 32086 26130
tri 31813 26119 31821 26127 ne
rect 31821 26122 32086 26127
tri 32086 26122 32094 26130 sw
rect 70802 26124 71000 26182
rect 31821 26119 32094 26122
tri 31821 26111 31829 26119 ne
rect 31829 26114 32094 26119
tri 32094 26114 32102 26122 sw
rect 31829 26111 32102 26114
tri 31829 26103 31837 26111 ne
rect 31837 26106 32102 26111
tri 32102 26106 32110 26114 sw
rect 31837 26103 32110 26106
tri 31837 26099 31841 26103 ne
rect 31841 26099 32110 26103
tri 31841 26091 31849 26099 ne
rect 31849 26098 32110 26099
tri 32110 26098 32118 26106 sw
rect 31849 26091 32118 26098
tri 31849 26083 31857 26091 ne
rect 31857 26090 32118 26091
tri 32118 26090 32126 26098 sw
rect 31857 26083 32126 26090
tri 31857 26075 31865 26083 ne
rect 31865 26082 32126 26083
tri 32126 26082 32134 26090 sw
rect 31865 26080 32134 26082
rect 31865 26075 31998 26080
tri 31865 26067 31873 26075 ne
rect 31873 26067 31998 26075
tri 31873 26059 31881 26067 ne
rect 31881 26059 31998 26067
tri 31881 26051 31889 26059 ne
rect 31889 26051 31998 26059
tri 31889 26043 31897 26051 ne
rect 31897 26043 31998 26051
tri 31897 26035 31905 26043 ne
rect 31905 26035 31998 26043
tri 31905 26027 31913 26035 ne
rect 31913 26034 31998 26035
rect 32044 26074 32134 26080
tri 32134 26074 32142 26082 sw
rect 70802 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26066 32142 26074
tri 32142 26066 32150 26074 sw
rect 32044 26058 32150 26066
tri 32150 26058 32158 26066 sw
rect 32044 26050 32158 26058
tri 32158 26050 32166 26058 sw
rect 32044 26042 32166 26050
tri 32166 26042 32174 26050 sw
rect 32044 26037 32174 26042
tri 32174 26037 32179 26042 sw
rect 32044 26034 32179 26037
rect 31913 26029 32179 26034
tri 32179 26029 32187 26037 sw
rect 31913 26027 32187 26029
tri 31913 26019 31921 26027 ne
rect 31921 26021 32187 26027
tri 32187 26021 32195 26029 sw
rect 31921 26019 32195 26021
tri 31921 26011 31929 26019 ne
rect 31929 26013 32195 26019
tri 32195 26013 32203 26021 sw
rect 70802 26020 71000 26078
rect 31929 26011 32203 26013
tri 31929 26003 31937 26011 ne
rect 31937 26005 32203 26011
tri 32203 26005 32211 26013 sw
rect 31937 26003 32211 26005
tri 31937 25995 31945 26003 ne
rect 31945 25997 32211 26003
tri 32211 25997 32219 26005 sw
rect 31945 25995 32219 25997
tri 31945 25987 31953 25995 ne
rect 31953 25989 32219 25995
tri 32219 25989 32227 25997 sw
rect 31953 25987 32227 25989
tri 31953 25979 31961 25987 ne
rect 31961 25981 32227 25987
tri 32227 25981 32235 25989 sw
rect 31961 25979 32235 25981
tri 31961 25971 31969 25979 ne
rect 31969 25973 32235 25979
tri 32235 25973 32243 25981 sw
rect 70802 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 31969 25971 32243 25973
tri 31969 25963 31977 25971 ne
rect 31977 25965 32243 25971
tri 32243 25965 32251 25973 sw
rect 31977 25963 32251 25965
tri 32251 25963 32253 25965 sw
tri 31977 25961 31979 25963 ne
rect 31979 25961 32253 25963
tri 31979 25955 31985 25961 ne
rect 31985 25955 32253 25961
tri 32253 25955 32261 25963 sw
tri 31985 25947 31993 25955 ne
rect 31993 25948 32261 25955
rect 31993 25947 32130 25948
tri 31993 25939 32001 25947 ne
rect 32001 25939 32130 25947
tri 32001 25931 32009 25939 ne
rect 32009 25931 32130 25939
tri 32009 25923 32017 25931 ne
rect 32017 25923 32130 25931
tri 32017 25915 32025 25923 ne
rect 32025 25915 32130 25923
tri 32025 25907 32033 25915 ne
rect 32033 25907 32130 25915
tri 32033 25899 32041 25907 ne
rect 32041 25902 32130 25907
rect 32176 25947 32261 25948
tri 32261 25947 32269 25955 sw
rect 32176 25939 32269 25947
tri 32269 25939 32277 25947 sw
rect 32176 25931 32277 25939
tri 32277 25931 32285 25939 sw
rect 32176 25923 32285 25931
tri 32285 25923 32293 25931 sw
rect 32176 25915 32293 25923
tri 32293 25915 32301 25923 sw
rect 70802 25916 71000 25974
rect 32176 25907 32301 25915
tri 32301 25907 32309 25915 sw
rect 32176 25902 32309 25907
rect 32041 25899 32309 25902
tri 32309 25899 32317 25907 sw
tri 32041 25894 32046 25899 ne
rect 32046 25894 32317 25899
tri 32046 25886 32054 25894 ne
rect 32054 25891 32317 25894
tri 32317 25891 32325 25899 sw
rect 32054 25886 32325 25891
tri 32325 25886 32330 25891 sw
tri 32054 25878 32062 25886 ne
rect 32062 25878 32330 25886
tri 32330 25878 32338 25886 sw
tri 32062 25870 32070 25878 ne
rect 32070 25870 32338 25878
tri 32338 25870 32346 25878 sw
rect 70802 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32070 25862 32078 25870 ne
rect 32078 25862 32346 25870
tri 32346 25862 32354 25870 sw
tri 32078 25854 32086 25862 ne
rect 32086 25854 32354 25862
tri 32354 25854 32362 25862 sw
tri 32086 25846 32094 25854 ne
rect 32094 25846 32362 25854
tri 32362 25846 32370 25854 sw
tri 32094 25838 32102 25846 ne
rect 32102 25838 32370 25846
tri 32370 25838 32378 25846 sw
tri 32102 25830 32110 25838 ne
rect 32110 25830 32378 25838
tri 32378 25830 32386 25838 sw
tri 32110 25822 32118 25830 ne
rect 32118 25822 32386 25830
tri 32386 25822 32394 25830 sw
tri 32118 25814 32126 25822 ne
rect 32126 25816 32394 25822
rect 32126 25814 32262 25816
tri 32126 25806 32134 25814 ne
rect 32134 25806 32262 25814
tri 32134 25798 32142 25806 ne
rect 32142 25798 32262 25806
tri 32142 25790 32150 25798 ne
rect 32150 25790 32262 25798
tri 32150 25782 32158 25790 ne
rect 32158 25782 32262 25790
tri 32158 25774 32166 25782 ne
rect 32166 25774 32262 25782
tri 32166 25766 32174 25774 ne
rect 32174 25770 32262 25774
rect 32308 25814 32394 25816
tri 32394 25814 32402 25822 sw
rect 32308 25806 32402 25814
tri 32402 25806 32410 25814 sw
rect 70802 25812 71000 25870
rect 32308 25798 32410 25806
tri 32410 25798 32418 25806 sw
rect 32308 25790 32418 25798
tri 32418 25790 32426 25798 sw
rect 32308 25782 32426 25790
tri 32426 25782 32434 25790 sw
rect 32308 25774 32434 25782
tri 32434 25774 32442 25782 sw
rect 32308 25771 32442 25774
tri 32442 25771 32445 25774 sw
rect 32308 25770 32445 25771
rect 32174 25766 32445 25770
tri 32174 25758 32182 25766 ne
rect 32182 25763 32445 25766
tri 32445 25763 32453 25771 sw
rect 70802 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 32182 25758 32453 25763
tri 32182 25750 32190 25758 ne
rect 32190 25755 32453 25758
tri 32453 25755 32461 25763 sw
rect 32190 25750 32461 25755
tri 32190 25742 32198 25750 ne
rect 32198 25747 32461 25750
tri 32461 25747 32469 25755 sw
rect 32198 25742 32469 25747
tri 32198 25734 32206 25742 ne
rect 32206 25739 32469 25742
tri 32469 25739 32477 25747 sw
rect 32206 25734 32477 25739
tri 32206 25726 32214 25734 ne
rect 32214 25731 32477 25734
tri 32477 25731 32485 25739 sw
rect 32214 25726 32485 25731
tri 32214 25718 32222 25726 ne
rect 32222 25723 32485 25726
tri 32485 25723 32493 25731 sw
rect 32222 25718 32493 25723
tri 32222 25711 32229 25718 ne
rect 32229 25715 32493 25718
tri 32493 25715 32501 25723 sw
rect 32229 25711 32501 25715
tri 32229 25703 32237 25711 ne
rect 32237 25707 32501 25711
tri 32501 25707 32509 25715 sw
rect 70802 25708 71000 25766
rect 32237 25703 32509 25707
tri 32509 25703 32513 25707 sw
tri 32237 25695 32245 25703 ne
rect 32245 25699 32513 25703
tri 32513 25699 32517 25703 sw
rect 32245 25695 32517 25699
tri 32245 25687 32253 25695 ne
rect 32253 25691 32517 25695
tri 32517 25691 32525 25699 sw
rect 32253 25687 32525 25691
tri 32253 25679 32261 25687 ne
rect 32261 25684 32525 25687
rect 32261 25679 32394 25684
tri 32261 25671 32269 25679 ne
rect 32269 25671 32394 25679
tri 32269 25663 32277 25671 ne
rect 32277 25663 32394 25671
tri 32277 25655 32285 25663 ne
rect 32285 25655 32394 25663
tri 32285 25647 32293 25655 ne
rect 32293 25647 32394 25655
tri 32293 25639 32301 25647 ne
rect 32301 25639 32394 25647
tri 32301 25631 32309 25639 ne
rect 32309 25638 32394 25639
rect 32440 25683 32525 25684
tri 32525 25683 32533 25691 sw
rect 32440 25675 32533 25683
tri 32533 25675 32541 25683 sw
rect 32440 25667 32541 25675
tri 32541 25667 32549 25675 sw
rect 32440 25659 32549 25667
tri 32549 25659 32557 25667 sw
rect 70802 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25651 32557 25659
tri 32557 25651 32565 25659 sw
rect 32440 25643 32565 25651
tri 32565 25643 32573 25651 sw
rect 32440 25638 32573 25643
rect 32309 25635 32573 25638
tri 32573 25635 32581 25643 sw
rect 32309 25634 32581 25635
tri 32581 25634 32582 25635 sw
rect 32309 25631 32582 25634
tri 32309 25626 32314 25631 ne
rect 32314 25626 32582 25631
tri 32582 25626 32590 25634 sw
tri 32314 25618 32322 25626 ne
rect 32322 25618 32590 25626
tri 32590 25618 32598 25626 sw
tri 32322 25610 32330 25618 ne
rect 32330 25610 32598 25618
tri 32598 25610 32606 25618 sw
tri 32330 25602 32338 25610 ne
rect 32338 25602 32606 25610
tri 32606 25602 32614 25610 sw
rect 70802 25604 71000 25662
tri 32338 25594 32346 25602 ne
rect 32346 25594 32614 25602
tri 32614 25594 32622 25602 sw
tri 32346 25586 32354 25594 ne
rect 32354 25586 32622 25594
tri 32622 25586 32630 25594 sw
tri 32354 25578 32362 25586 ne
rect 32362 25578 32630 25586
tri 32630 25578 32638 25586 sw
tri 32362 25570 32370 25578 ne
rect 32370 25570 32638 25578
tri 32638 25570 32646 25578 sw
tri 32370 25562 32378 25570 ne
rect 32378 25562 32646 25570
tri 32646 25562 32654 25570 sw
tri 32378 25554 32386 25562 ne
rect 32386 25554 32654 25562
tri 32654 25554 32662 25562 sw
rect 70802 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
tri 32386 25546 32394 25554 ne
rect 32394 25552 32662 25554
rect 32394 25546 32526 25552
tri 32394 25538 32402 25546 ne
rect 32402 25538 32526 25546
tri 32402 25530 32410 25538 ne
rect 32410 25530 32526 25538
tri 32410 25522 32418 25530 ne
rect 32418 25522 32526 25530
tri 32418 25514 32426 25522 ne
rect 32426 25514 32526 25522
tri 32426 25506 32434 25514 ne
rect 32434 25506 32526 25514
rect 32572 25546 32662 25552
tri 32662 25546 32670 25554 sw
rect 32572 25538 32670 25546
tri 32670 25538 32678 25546 sw
rect 32572 25530 32678 25538
tri 32678 25530 32686 25538 sw
rect 32572 25522 32686 25530
tri 32686 25522 32694 25530 sw
rect 32572 25514 32694 25522
tri 32694 25514 32702 25522 sw
rect 32572 25512 32702 25514
tri 32702 25512 32704 25514 sw
rect 32572 25506 32704 25512
tri 32434 25499 32441 25506 ne
rect 32441 25504 32704 25506
tri 32704 25504 32712 25512 sw
rect 32441 25499 32712 25504
tri 32441 25491 32449 25499 ne
rect 32449 25496 32712 25499
tri 32712 25496 32720 25504 sw
rect 70802 25500 71000 25558
rect 32449 25491 32720 25496
tri 32449 25483 32457 25491 ne
rect 32457 25488 32720 25491
tri 32720 25488 32728 25496 sw
rect 32457 25483 32728 25488
tri 32457 25475 32465 25483 ne
rect 32465 25480 32728 25483
tri 32728 25480 32736 25488 sw
rect 32465 25475 32736 25480
tri 32465 25467 32473 25475 ne
rect 32473 25472 32736 25475
tri 32736 25472 32744 25480 sw
rect 32473 25467 32744 25472
tri 32473 25459 32481 25467 ne
rect 32481 25464 32744 25467
tri 32744 25464 32752 25472 sw
rect 32481 25459 32752 25464
tri 32481 25451 32489 25459 ne
rect 32489 25456 32752 25459
tri 32752 25456 32760 25464 sw
rect 32489 25451 32760 25456
tri 32489 25443 32497 25451 ne
rect 32497 25448 32760 25451
tri 32760 25448 32768 25456 sw
rect 70802 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32497 25443 32768 25448
tri 32497 25435 32505 25443 ne
rect 32505 25440 32768 25443
tri 32768 25440 32776 25448 sw
rect 32505 25439 32776 25440
tri 32776 25439 32777 25440 sw
rect 32505 25435 32777 25439
tri 32505 25431 32509 25435 ne
rect 32509 25431 32777 25435
tri 32777 25431 32785 25439 sw
tri 32509 25423 32517 25431 ne
rect 32517 25423 32785 25431
tri 32785 25423 32793 25431 sw
tri 32517 25415 32525 25423 ne
rect 32525 25420 32793 25423
rect 32525 25415 32658 25420
tri 32525 25407 32533 25415 ne
rect 32533 25407 32658 25415
tri 32533 25399 32541 25407 ne
rect 32541 25399 32658 25407
tri 32541 25391 32549 25399 ne
rect 32549 25391 32658 25399
tri 32549 25383 32557 25391 ne
rect 32557 25383 32658 25391
tri 32557 25375 32565 25383 ne
rect 32565 25375 32658 25383
tri 32565 25367 32573 25375 ne
rect 32573 25374 32658 25375
rect 32704 25415 32793 25420
tri 32793 25415 32801 25423 sw
rect 32704 25407 32801 25415
tri 32801 25407 32809 25415 sw
rect 32704 25399 32809 25407
tri 32809 25399 32817 25407 sw
rect 32704 25391 32817 25399
tri 32817 25391 32825 25399 sw
rect 70802 25396 71000 25454
rect 32704 25383 32825 25391
tri 32825 25383 32833 25391 sw
rect 32704 25375 32833 25383
tri 32833 25375 32841 25383 sw
rect 32704 25374 32841 25375
rect 32573 25371 32841 25374
tri 32841 25371 32845 25375 sw
rect 32573 25367 32845 25371
tri 32573 25359 32581 25367 ne
rect 32581 25363 32845 25367
tri 32845 25363 32853 25371 sw
rect 32581 25359 32853 25363
tri 32581 25351 32589 25359 ne
rect 32589 25355 32853 25359
tri 32853 25355 32861 25363 sw
rect 32589 25351 32861 25355
tri 32589 25346 32594 25351 ne
rect 32594 25347 32861 25351
tri 32861 25347 32869 25355 sw
rect 70802 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
rect 32594 25346 32869 25347
tri 32594 25338 32602 25346 ne
rect 32602 25339 32869 25346
tri 32869 25339 32877 25347 sw
rect 32602 25338 32877 25339
tri 32602 25330 32610 25338 ne
rect 32610 25331 32877 25338
tri 32877 25331 32885 25339 sw
rect 32610 25330 32885 25331
tri 32610 25322 32618 25330 ne
rect 32618 25323 32885 25330
tri 32885 25323 32893 25331 sw
rect 32618 25322 32893 25323
tri 32618 25314 32626 25322 ne
rect 32626 25315 32893 25322
tri 32893 25315 32901 25323 sw
rect 32626 25314 32901 25315
tri 32626 25306 32634 25314 ne
rect 32634 25307 32901 25314
tri 32901 25307 32909 25315 sw
rect 32634 25306 32909 25307
tri 32634 25298 32642 25306 ne
rect 32642 25299 32909 25306
tri 32909 25299 32917 25307 sw
rect 32642 25298 32917 25299
tri 32642 25290 32650 25298 ne
rect 32650 25291 32917 25298
tri 32917 25291 32925 25299 sw
rect 70802 25292 71000 25350
rect 32650 25290 32925 25291
tri 32650 25282 32658 25290 ne
rect 32658 25288 32925 25290
rect 32658 25282 32790 25288
tri 32658 25274 32666 25282 ne
rect 32666 25274 32790 25282
tri 32666 25266 32674 25274 ne
rect 32674 25266 32790 25274
tri 32674 25258 32682 25266 ne
rect 32682 25258 32790 25266
tri 32682 25250 32690 25258 ne
rect 32690 25250 32790 25258
tri 32690 25242 32698 25250 ne
rect 32698 25242 32790 25250
rect 32836 25283 32925 25288
tri 32925 25283 32933 25291 sw
rect 32836 25275 32933 25283
tri 32933 25275 32941 25283 sw
rect 32836 25267 32941 25275
tri 32941 25267 32949 25275 sw
rect 32836 25260 32949 25267
tri 32949 25260 32956 25267 sw
rect 32836 25252 32956 25260
tri 32956 25252 32964 25260 sw
rect 32836 25244 32964 25252
tri 32964 25244 32972 25252 sw
rect 70802 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 32836 25242 32972 25244
tri 32698 25234 32706 25242 ne
rect 32706 25236 32972 25242
tri 32972 25236 32980 25244 sw
rect 32706 25234 32980 25236
tri 32706 25226 32714 25234 ne
rect 32714 25228 32980 25234
tri 32980 25228 32988 25236 sw
rect 32714 25226 32988 25228
tri 32714 25218 32722 25226 ne
rect 32722 25220 32988 25226
tri 32988 25220 32996 25228 sw
rect 32722 25218 32996 25220
tri 32722 25215 32725 25218 ne
rect 32725 25215 32996 25218
tri 32725 25207 32733 25215 ne
rect 32733 25212 32996 25215
tri 32996 25212 33004 25220 sw
rect 32733 25207 33004 25212
tri 32733 25199 32741 25207 ne
rect 32741 25204 33004 25207
tri 33004 25204 33012 25212 sw
rect 32741 25199 33012 25204
tri 32741 25191 32749 25199 ne
rect 32749 25196 33012 25199
tri 33012 25196 33020 25204 sw
rect 32749 25191 33020 25196
tri 32749 25183 32757 25191 ne
rect 32757 25188 33020 25191
tri 33020 25188 33028 25196 sw
rect 70802 25188 71000 25246
rect 32757 25183 33028 25188
tri 32757 25175 32765 25183 ne
rect 32765 25180 33028 25183
tri 33028 25180 33036 25188 sw
rect 32765 25175 33036 25180
tri 32765 25167 32773 25175 ne
rect 32773 25172 33036 25175
tri 33036 25172 33044 25180 sw
rect 32773 25167 33044 25172
tri 32773 25159 32781 25167 ne
rect 32781 25164 33044 25167
tri 33044 25164 33052 25172 sw
rect 32781 25159 33052 25164
tri 32781 25151 32789 25159 ne
rect 32789 25156 33052 25159
tri 33052 25156 33060 25164 sw
rect 32789 25151 32922 25156
tri 32789 25143 32797 25151 ne
rect 32797 25143 32922 25151
tri 32797 25139 32801 25143 ne
rect 32801 25139 32922 25143
tri 32801 25131 32809 25139 ne
rect 32809 25131 32922 25139
tri 32809 25123 32817 25131 ne
rect 32817 25123 32922 25131
tri 32817 25115 32825 25123 ne
rect 32825 25115 32922 25123
tri 32825 25107 32833 25115 ne
rect 32833 25110 32922 25115
rect 32968 25155 33060 25156
tri 33060 25155 33061 25156 sw
rect 32968 25147 33061 25155
tri 33061 25147 33069 25155 sw
rect 32968 25139 33069 25147
tri 33069 25139 33077 25147 sw
rect 70802 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 32968 25131 33077 25139
tri 33077 25131 33085 25139 sw
rect 32968 25123 33085 25131
tri 33085 25123 33093 25131 sw
rect 32968 25115 33093 25123
tri 33093 25115 33101 25123 sw
rect 32968 25110 33101 25115
rect 32833 25107 33101 25110
tri 33101 25107 33109 25115 sw
tri 32833 25099 32841 25107 ne
rect 32841 25099 33109 25107
tri 33109 25099 33117 25107 sw
tri 32841 25091 32849 25099 ne
rect 32849 25091 33117 25099
tri 33117 25091 33125 25099 sw
tri 32849 25083 32857 25091 ne
rect 32857 25083 33125 25091
tri 33125 25083 33133 25091 sw
rect 70802 25084 71000 25142
tri 32857 25075 32865 25083 ne
rect 32865 25075 33133 25083
tri 33133 25075 33141 25083 sw
tri 32865 25067 32873 25075 ne
rect 32873 25067 33141 25075
tri 33141 25067 33149 25075 sw
tri 32873 25059 32881 25067 ne
rect 32881 25059 33149 25067
tri 33149 25059 33157 25067 sw
tri 32881 25051 32889 25059 ne
rect 32889 25051 33157 25059
tri 33157 25051 33165 25059 sw
tri 32889 25043 32897 25051 ne
rect 32897 25043 33165 25051
tri 33165 25043 33173 25051 sw
tri 32897 25035 32905 25043 ne
rect 32905 25035 33173 25043
tri 33173 25035 33181 25043 sw
rect 70802 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
tri 32905 25027 32913 25035 ne
rect 32913 25027 33181 25035
tri 33181 25027 33189 25035 sw
tri 32913 25019 32921 25027 ne
rect 32921 25024 33189 25027
rect 32921 25019 33054 25024
tri 32921 25016 32924 25019 ne
rect 32924 25016 33054 25019
tri 32924 25008 32932 25016 ne
rect 32932 25008 33054 25016
tri 32932 25000 32940 25008 ne
rect 32940 25000 33054 25008
tri 32940 24992 32948 25000 ne
rect 32948 24992 33054 25000
tri 32948 24984 32956 24992 ne
rect 32956 24984 33054 24992
tri 32956 24976 32964 24984 ne
rect 32964 24978 33054 24984
rect 33100 25019 33189 25024
tri 33189 25019 33197 25027 sw
rect 33100 25016 33197 25019
tri 33197 25016 33200 25019 sw
rect 33100 25008 33200 25016
tri 33200 25008 33208 25016 sw
rect 33100 25000 33208 25008
tri 33208 25000 33216 25008 sw
rect 33100 24992 33216 25000
tri 33216 24992 33224 25000 sw
rect 33100 24984 33224 24992
tri 33224 24984 33232 24992 sw
rect 33100 24978 33232 24984
rect 32964 24976 33232 24978
tri 33232 24976 33240 24984 sw
rect 70802 24980 71000 25038
tri 32964 24968 32972 24976 ne
rect 32972 24968 33240 24976
tri 33240 24968 33248 24976 sw
tri 32972 24960 32980 24968 ne
rect 32980 24960 33248 24968
tri 33248 24960 33256 24968 sw
tri 32980 24952 32988 24960 ne
rect 32988 24952 33256 24960
tri 33256 24952 33264 24960 sw
tri 32988 24944 32996 24952 ne
rect 32996 24944 33264 24952
tri 33264 24944 33272 24952 sw
tri 32996 24936 33004 24944 ne
rect 33004 24936 33272 24944
tri 33272 24936 33280 24944 sw
tri 33004 24928 33012 24936 ne
rect 33012 24928 33280 24936
tri 33280 24928 33288 24936 sw
rect 70802 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33012 24920 33020 24928 ne
rect 33020 24920 33288 24928
tri 33288 24920 33296 24928 sw
tri 33020 24912 33028 24920 ne
rect 33028 24912 33296 24920
tri 33296 24912 33304 24920 sw
tri 33028 24911 33029 24912 ne
rect 33029 24911 33304 24912
tri 33304 24911 33305 24912 sw
tri 33029 24903 33037 24911 ne
rect 33037 24903 33305 24911
tri 33305 24903 33313 24911 sw
tri 33037 24895 33045 24903 ne
rect 33045 24895 33313 24903
tri 33313 24895 33321 24903 sw
tri 33045 24887 33053 24895 ne
rect 33053 24892 33321 24895
rect 33053 24887 33186 24892
tri 33053 24879 33061 24887 ne
rect 33061 24879 33186 24887
tri 33061 24871 33069 24879 ne
rect 33069 24871 33186 24879
tri 33069 24863 33077 24871 ne
rect 33077 24863 33186 24871
tri 33077 24855 33085 24863 ne
rect 33085 24855 33186 24863
tri 33085 24847 33093 24855 ne
rect 33093 24847 33186 24855
tri 33093 24839 33101 24847 ne
rect 33101 24846 33186 24847
rect 33232 24887 33321 24892
tri 33321 24887 33329 24895 sw
rect 33232 24879 33329 24887
tri 33329 24879 33337 24887 sw
rect 33232 24871 33337 24879
tri 33337 24871 33345 24879 sw
rect 70802 24876 71000 24934
rect 33232 24863 33345 24871
tri 33345 24863 33353 24871 sw
rect 33232 24855 33353 24863
tri 33353 24855 33361 24863 sw
rect 33232 24847 33361 24855
tri 33361 24847 33369 24855 sw
rect 33232 24846 33369 24847
rect 33101 24839 33369 24846
tri 33369 24839 33377 24847 sw
tri 33101 24831 33109 24839 ne
rect 33109 24833 33377 24839
tri 33377 24833 33383 24839 sw
rect 33109 24831 33383 24833
tri 33109 24823 33117 24831 ne
rect 33117 24825 33383 24831
tri 33383 24825 33391 24833 sw
rect 70802 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 33117 24823 33391 24825
tri 33117 24818 33122 24823 ne
rect 33122 24818 33391 24823
tri 33122 24810 33130 24818 ne
rect 33130 24817 33391 24818
tri 33391 24817 33399 24825 sw
rect 33130 24810 33399 24817
tri 33130 24802 33138 24810 ne
rect 33138 24809 33399 24810
tri 33399 24809 33407 24817 sw
rect 33138 24802 33407 24809
tri 33138 24794 33146 24802 ne
rect 33146 24801 33407 24802
tri 33407 24801 33415 24809 sw
rect 33146 24794 33415 24801
tri 33146 24786 33154 24794 ne
rect 33154 24793 33415 24794
tri 33415 24793 33423 24801 sw
rect 33154 24786 33423 24793
tri 33154 24778 33162 24786 ne
rect 33162 24785 33423 24786
tri 33423 24785 33431 24793 sw
rect 33162 24778 33431 24785
tri 33162 24770 33170 24778 ne
rect 33170 24777 33431 24778
tri 33431 24777 33439 24785 sw
rect 33170 24770 33439 24777
tri 33170 24762 33178 24770 ne
rect 33178 24769 33439 24770
tri 33439 24769 33447 24777 sw
rect 70802 24772 71000 24830
rect 33178 24762 33447 24769
tri 33178 24754 33186 24762 ne
rect 33186 24761 33447 24762
tri 33447 24761 33455 24769 sw
rect 33186 24760 33455 24761
rect 33186 24754 33318 24760
tri 33186 24746 33194 24754 ne
rect 33194 24746 33318 24754
tri 33194 24738 33202 24746 ne
rect 33202 24738 33318 24746
tri 33202 24730 33210 24738 ne
rect 33210 24730 33318 24738
tri 33210 24722 33218 24730 ne
rect 33218 24722 33318 24730
tri 33218 24714 33226 24722 ne
rect 33226 24714 33318 24722
rect 33364 24753 33455 24760
tri 33455 24753 33463 24761 sw
rect 33364 24745 33463 24753
tri 33463 24745 33471 24753 sw
rect 33364 24737 33471 24745
tri 33471 24737 33479 24745 sw
rect 33364 24729 33479 24737
tri 33479 24729 33487 24737 sw
rect 33364 24721 33487 24729
tri 33487 24721 33495 24729 sw
rect 70802 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 33364 24714 33495 24721
tri 33226 24706 33234 24714 ne
rect 33234 24713 33495 24714
tri 33495 24713 33503 24721 sw
rect 33234 24708 33503 24713
tri 33503 24708 33508 24713 sw
rect 33234 24706 33508 24708
tri 33234 24698 33242 24706 ne
rect 33242 24700 33508 24706
tri 33508 24700 33516 24708 sw
rect 33242 24698 33516 24700
tri 33242 24690 33250 24698 ne
rect 33250 24692 33516 24698
tri 33516 24692 33524 24700 sw
rect 33250 24690 33524 24692
tri 33250 24688 33252 24690 ne
rect 33252 24688 33524 24690
tri 33252 24680 33260 24688 ne
rect 33260 24684 33524 24688
tri 33524 24684 33532 24692 sw
rect 33260 24680 33532 24684
tri 33260 24672 33268 24680 ne
rect 33268 24676 33532 24680
tri 33532 24676 33540 24684 sw
rect 33268 24672 33540 24676
tri 33268 24664 33276 24672 ne
rect 33276 24668 33540 24672
tri 33540 24668 33548 24676 sw
rect 70802 24668 71000 24726
rect 33276 24664 33548 24668
tri 33276 24656 33284 24664 ne
rect 33284 24660 33548 24664
tri 33548 24660 33556 24668 sw
rect 33284 24656 33556 24660
tri 33284 24648 33292 24656 ne
rect 33292 24652 33556 24656
tri 33556 24652 33564 24660 sw
rect 33292 24648 33564 24652
tri 33292 24640 33300 24648 ne
rect 33300 24644 33564 24648
tri 33564 24644 33572 24652 sw
rect 33300 24640 33572 24644
tri 33300 24632 33308 24640 ne
rect 33308 24636 33572 24640
tri 33572 24636 33580 24644 sw
rect 33308 24632 33580 24636
tri 33308 24624 33316 24632 ne
rect 33316 24628 33580 24632
tri 33580 24628 33588 24636 sw
rect 33316 24624 33450 24628
tri 33316 24619 33321 24624 ne
rect 33321 24619 33450 24624
tri 33321 24611 33329 24619 ne
rect 33329 24611 33450 24619
tri 33329 24603 33337 24611 ne
rect 33337 24603 33450 24611
tri 33337 24595 33345 24603 ne
rect 33345 24595 33450 24603
tri 33345 24587 33353 24595 ne
rect 33353 24587 33450 24595
tri 33353 24579 33361 24587 ne
rect 33361 24582 33450 24587
rect 33496 24627 33588 24628
tri 33588 24627 33589 24628 sw
rect 33496 24619 33589 24627
tri 33589 24619 33597 24627 sw
rect 70802 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24611 33597 24619
tri 33597 24611 33605 24619 sw
rect 33496 24603 33605 24611
tri 33605 24603 33613 24611 sw
rect 33496 24595 33613 24603
tri 33613 24595 33621 24603 sw
rect 33496 24587 33621 24595
tri 33621 24587 33629 24595 sw
rect 33496 24582 33629 24587
rect 33361 24579 33629 24582
tri 33629 24579 33637 24587 sw
tri 33361 24571 33369 24579 ne
rect 33369 24571 33637 24579
tri 33637 24571 33645 24579 sw
tri 33369 24563 33377 24571 ne
rect 33377 24563 33645 24571
tri 33645 24563 33653 24571 sw
rect 70802 24564 71000 24622
tri 33377 24555 33385 24563 ne
rect 33385 24555 33653 24563
tri 33653 24555 33661 24563 sw
tri 33385 24547 33393 24555 ne
rect 33393 24551 33661 24555
tri 33661 24551 33665 24555 sw
rect 33393 24547 33665 24551
tri 33393 24546 33394 24547 ne
rect 33394 24546 33665 24547
tri 33394 24538 33402 24546 ne
rect 33402 24543 33665 24546
tri 33665 24543 33673 24551 sw
rect 33402 24538 33673 24543
tri 33402 24530 33410 24538 ne
rect 33410 24535 33673 24538
tri 33673 24535 33681 24543 sw
rect 33410 24530 33681 24535
tri 33410 24522 33418 24530 ne
rect 33418 24527 33681 24530
tri 33681 24527 33689 24535 sw
rect 33418 24522 33689 24527
tri 33418 24514 33426 24522 ne
rect 33426 24519 33689 24522
tri 33689 24519 33697 24527 sw
rect 33426 24514 33697 24519
tri 33426 24506 33434 24514 ne
rect 33434 24511 33697 24514
tri 33697 24511 33705 24519 sw
rect 70802 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
rect 33434 24506 33705 24511
tri 33434 24498 33442 24506 ne
rect 33442 24503 33705 24506
tri 33705 24503 33713 24511 sw
rect 33442 24498 33713 24503
tri 33442 24490 33450 24498 ne
rect 33450 24496 33713 24498
rect 33450 24490 33582 24496
tri 33450 24482 33458 24490 ne
rect 33458 24482 33582 24490
tri 33458 24474 33466 24482 ne
rect 33466 24474 33582 24482
tri 33466 24466 33474 24474 ne
rect 33474 24466 33582 24474
tri 33474 24458 33482 24466 ne
rect 33482 24458 33582 24466
tri 33482 24450 33490 24458 ne
rect 33490 24450 33582 24458
rect 33628 24495 33713 24496
tri 33713 24495 33721 24503 sw
rect 33628 24487 33721 24495
tri 33721 24487 33729 24495 sw
rect 33628 24479 33729 24487
tri 33729 24479 33737 24487 sw
rect 33628 24471 33737 24479
tri 33737 24471 33745 24479 sw
rect 33628 24463 33745 24471
tri 33745 24463 33753 24471 sw
rect 33628 24455 33753 24463
tri 33753 24455 33761 24463 sw
rect 70802 24460 71000 24518
rect 33628 24450 33761 24455
tri 33490 24442 33498 24450 ne
rect 33498 24447 33761 24450
tri 33761 24447 33769 24455 sw
rect 33498 24442 33769 24447
tri 33498 24434 33506 24442 ne
rect 33506 24439 33769 24442
tri 33769 24439 33777 24447 sw
rect 33506 24434 33777 24439
tri 33777 24434 33782 24439 sw
tri 33506 24426 33514 24434 ne
rect 33514 24426 33782 24434
tri 33782 24426 33790 24434 sw
tri 33514 24418 33522 24426 ne
rect 33522 24418 33790 24426
tri 33790 24418 33798 24426 sw
tri 33522 24410 33530 24418 ne
rect 33530 24410 33798 24418
tri 33798 24410 33806 24418 sw
rect 70802 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33530 24402 33538 24410 ne
rect 33538 24402 33806 24410
tri 33806 24402 33814 24410 sw
tri 33538 24394 33546 24402 ne
rect 33546 24394 33814 24402
tri 33814 24394 33822 24402 sw
tri 33546 24386 33554 24394 ne
rect 33554 24386 33822 24394
tri 33822 24386 33830 24394 sw
tri 33554 24378 33562 24386 ne
rect 33562 24378 33830 24386
tri 33830 24378 33838 24386 sw
tri 33562 24370 33570 24378 ne
rect 33570 24370 33838 24378
tri 33838 24370 33846 24378 sw
tri 33570 24366 33574 24370 ne
rect 33574 24366 33846 24370
tri 33846 24366 33850 24370 sw
tri 33574 24362 33578 24366 ne
rect 33578 24364 33850 24366
rect 33578 24362 33714 24364
tri 33578 24354 33586 24362 ne
rect 33586 24354 33714 24362
tri 33586 24346 33594 24354 ne
rect 33594 24346 33714 24354
tri 33594 24338 33602 24346 ne
rect 33602 24338 33714 24346
tri 33602 24330 33610 24338 ne
rect 33610 24330 33714 24338
tri 33610 24322 33618 24330 ne
rect 33618 24322 33714 24330
tri 33618 24314 33626 24322 ne
rect 33626 24318 33714 24322
rect 33760 24362 33850 24364
tri 33850 24362 33854 24366 sw
rect 33760 24354 33854 24362
tri 33854 24354 33862 24362 sw
rect 70802 24356 71000 24414
rect 33760 24346 33862 24354
tri 33862 24346 33870 24354 sw
rect 33760 24338 33870 24346
tri 33870 24338 33878 24346 sw
rect 33760 24330 33878 24338
tri 33878 24330 33886 24338 sw
rect 33760 24322 33886 24330
tri 33886 24322 33894 24330 sw
rect 33760 24318 33894 24322
rect 33626 24314 33894 24318
tri 33894 24314 33902 24322 sw
tri 33626 24306 33634 24314 ne
rect 33634 24306 33902 24314
tri 33902 24306 33910 24314 sw
rect 70802 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
tri 33634 24298 33642 24306 ne
rect 33642 24298 33910 24306
tri 33910 24298 33918 24306 sw
tri 33642 24290 33650 24298 ne
rect 33650 24290 33918 24298
tri 33918 24290 33926 24298 sw
tri 33650 24282 33658 24290 ne
rect 33658 24282 33926 24290
tri 33926 24282 33934 24290 sw
tri 33658 24274 33666 24282 ne
rect 33666 24274 33934 24282
tri 33934 24274 33942 24282 sw
tri 33666 24266 33674 24274 ne
rect 33674 24266 33942 24274
tri 33942 24266 33950 24274 sw
tri 33674 24258 33682 24266 ne
rect 33682 24258 33950 24266
tri 33950 24258 33958 24266 sw
tri 33682 24250 33690 24258 ne
rect 33690 24250 33958 24258
tri 33958 24250 33966 24258 sw
rect 70802 24252 71000 24310
tri 33690 24249 33691 24250 ne
rect 33691 24249 33966 24250
tri 33966 24249 33967 24250 sw
tri 33691 24241 33699 24249 ne
rect 33699 24241 33967 24249
tri 33967 24241 33975 24249 sw
tri 33699 24233 33707 24241 ne
rect 33707 24233 33975 24241
tri 33975 24233 33983 24241 sw
tri 33707 24225 33715 24233 ne
rect 33715 24232 33983 24233
rect 33715 24225 33846 24232
tri 33715 24217 33723 24225 ne
rect 33723 24217 33846 24225
tri 33723 24209 33731 24217 ne
rect 33731 24209 33846 24217
tri 33731 24201 33739 24209 ne
rect 33739 24201 33846 24209
tri 33739 24193 33747 24201 ne
rect 33747 24193 33846 24201
tri 33747 24185 33755 24193 ne
rect 33755 24186 33846 24193
rect 33892 24225 33983 24232
tri 33983 24225 33991 24233 sw
rect 33892 24217 33991 24225
tri 33991 24217 33999 24225 sw
rect 33892 24209 33999 24217
tri 33999 24209 34007 24217 sw
rect 33892 24201 34007 24209
tri 34007 24201 34015 24209 sw
rect 70802 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 33892 24193 34015 24201
tri 34015 24193 34023 24201 sw
rect 33892 24186 34023 24193
rect 33755 24185 34023 24186
tri 34023 24185 34031 24193 sw
tri 33755 24177 33763 24185 ne
rect 33763 24177 34031 24185
tri 34031 24177 34039 24185 sw
tri 33763 24169 33771 24177 ne
rect 33771 24169 34039 24177
tri 34039 24169 34047 24177 sw
tri 33771 24161 33779 24169 ne
rect 33779 24161 34047 24169
tri 34047 24161 34055 24169 sw
tri 33779 24153 33787 24161 ne
rect 33787 24153 34055 24161
tri 34055 24153 34063 24161 sw
tri 33787 24145 33795 24153 ne
rect 33795 24145 34063 24153
tri 34063 24145 34071 24153 sw
rect 70802 24148 71000 24206
tri 33795 24137 33803 24145 ne
rect 33803 24137 34071 24145
tri 34071 24137 34079 24145 sw
tri 33803 24129 33811 24137 ne
rect 33811 24129 34079 24137
tri 34079 24129 34087 24137 sw
tri 33811 24121 33819 24129 ne
rect 33819 24121 34087 24129
tri 34087 24121 34095 24129 sw
tri 33819 24113 33827 24121 ne
rect 33827 24113 34095 24121
tri 34095 24113 34103 24121 sw
tri 33827 24107 33833 24113 ne
rect 33833 24107 34103 24113
tri 34103 24107 34109 24113 sw
tri 33833 24099 33841 24107 ne
rect 33841 24100 34109 24107
rect 33841 24099 33978 24100
tri 33841 24091 33849 24099 ne
rect 33849 24091 33978 24099
tri 33849 24086 33854 24091 ne
rect 33854 24086 33978 24091
tri 33854 24083 33857 24086 ne
rect 33857 24083 33978 24086
tri 33857 24075 33865 24083 ne
rect 33865 24075 33978 24083
tri 33865 24067 33873 24075 ne
rect 33873 24067 33978 24075
tri 33873 24059 33881 24067 ne
rect 33881 24059 33978 24067
tri 33881 24051 33889 24059 ne
rect 33889 24054 33978 24059
rect 34024 24099 34109 24100
tri 34109 24099 34117 24107 sw
rect 70802 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 34024 24091 34117 24099
tri 34117 24091 34125 24099 sw
rect 34024 24083 34125 24091
tri 34125 24083 34133 24091 sw
rect 34024 24075 34133 24083
tri 34133 24075 34141 24083 sw
rect 34024 24067 34141 24075
tri 34141 24067 34149 24075 sw
rect 34024 24059 34149 24067
tri 34149 24059 34157 24067 sw
rect 34024 24054 34157 24059
rect 33889 24051 34157 24054
tri 34157 24051 34165 24059 sw
tri 33889 24043 33897 24051 ne
rect 33897 24043 34165 24051
tri 34165 24043 34173 24051 sw
rect 70802 24044 71000 24102
tri 33897 24035 33905 24043 ne
rect 33905 24035 34173 24043
tri 34173 24035 34181 24043 sw
tri 33905 24027 33913 24035 ne
rect 33913 24027 34181 24035
tri 34181 24027 34189 24035 sw
tri 33913 24019 33921 24027 ne
rect 33921 24019 34189 24027
tri 34189 24019 34197 24027 sw
tri 33921 24011 33929 24019 ne
rect 33929 24011 34197 24019
tri 34197 24011 34205 24019 sw
tri 33929 24003 33937 24011 ne
rect 33937 24003 34205 24011
tri 34205 24003 34213 24011 sw
tri 33937 23995 33945 24003 ne
rect 33945 23995 34213 24003
tri 34213 23995 34221 24003 sw
rect 70802 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33945 23987 33953 23995 ne
rect 33953 23987 34221 23995
tri 34221 23987 34229 23995 sw
tri 33953 23979 33961 23987 ne
rect 33961 23979 34229 23987
tri 34229 23979 34237 23987 sw
tri 33961 23971 33969 23979 ne
rect 33969 23971 34237 23979
tri 34237 23971 34245 23979 sw
tri 33969 23967 33973 23971 ne
rect 33973 23968 34245 23971
rect 33973 23967 34110 23968
tri 33973 23959 33981 23967 ne
rect 33981 23959 34110 23967
tri 33981 23951 33989 23959 ne
rect 33989 23951 34110 23959
tri 33989 23943 33997 23951 ne
rect 33997 23943 34110 23951
tri 33997 23935 34005 23943 ne
rect 34005 23935 34110 23943
tri 34005 23927 34013 23935 ne
rect 34013 23927 34110 23935
tri 34013 23919 34021 23927 ne
rect 34021 23922 34110 23927
rect 34156 23965 34245 23968
tri 34245 23965 34251 23971 sw
rect 34156 23957 34251 23965
tri 34251 23957 34259 23965 sw
rect 34156 23949 34259 23957
tri 34259 23949 34267 23957 sw
rect 34156 23941 34267 23949
tri 34267 23941 34275 23949 sw
rect 34156 23933 34275 23941
tri 34275 23933 34283 23941 sw
rect 70802 23940 71000 23998
rect 34156 23925 34283 23933
tri 34283 23925 34291 23933 sw
rect 34156 23922 34291 23925
rect 34021 23919 34291 23922
tri 34021 23911 34029 23919 ne
rect 34029 23917 34291 23919
tri 34291 23917 34299 23925 sw
rect 34029 23911 34299 23917
tri 34029 23903 34037 23911 ne
rect 34037 23909 34299 23911
tri 34299 23909 34307 23917 sw
rect 34037 23903 34307 23909
tri 34037 23895 34045 23903 ne
rect 34045 23901 34307 23903
tri 34307 23901 34315 23909 sw
rect 34045 23895 34315 23901
tri 34045 23887 34053 23895 ne
rect 34053 23893 34315 23895
tri 34315 23893 34323 23901 sw
rect 70802 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
rect 34053 23887 34323 23893
tri 34053 23879 34061 23887 ne
rect 34061 23885 34323 23887
tri 34323 23885 34331 23893 sw
rect 34061 23879 34331 23885
tri 34061 23871 34069 23879 ne
rect 34069 23877 34331 23879
tri 34331 23877 34339 23885 sw
rect 34069 23871 34339 23877
tri 34069 23863 34077 23871 ne
rect 34077 23869 34339 23871
tri 34339 23869 34347 23877 sw
rect 34077 23863 34347 23869
tri 34077 23861 34079 23863 ne
rect 34079 23861 34347 23863
tri 34347 23861 34355 23869 sw
tri 34079 23855 34085 23861 ne
rect 34085 23855 34355 23861
tri 34355 23855 34361 23861 sw
tri 34085 23847 34093 23855 ne
rect 34093 23847 34361 23855
tri 34361 23847 34369 23855 sw
tri 34093 23839 34101 23847 ne
rect 34101 23839 34369 23847
tri 34369 23839 34377 23847 sw
tri 34101 23831 34109 23839 ne
rect 34109 23836 34377 23839
rect 34109 23831 34242 23836
tri 34109 23823 34117 23831 ne
rect 34117 23823 34242 23831
tri 34117 23815 34125 23823 ne
rect 34125 23815 34242 23823
tri 34125 23807 34133 23815 ne
rect 34133 23807 34242 23815
tri 34133 23799 34141 23807 ne
rect 34141 23799 34242 23807
tri 34141 23791 34149 23799 ne
rect 34149 23791 34242 23799
tri 34149 23783 34157 23791 ne
rect 34157 23790 34242 23791
rect 34288 23831 34377 23836
tri 34377 23831 34385 23839 sw
rect 70802 23836 71000 23894
rect 34288 23823 34385 23831
tri 34385 23823 34393 23831 sw
rect 34288 23815 34393 23823
tri 34393 23815 34401 23823 sw
rect 34288 23807 34401 23815
tri 34401 23807 34409 23815 sw
rect 34288 23799 34409 23807
tri 34409 23799 34417 23807 sw
rect 34288 23791 34417 23799
tri 34417 23791 34425 23799 sw
rect 34288 23790 34425 23791
rect 34157 23788 34425 23790
tri 34425 23788 34428 23791 sw
rect 70802 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
rect 34157 23783 34428 23788
tri 34157 23775 34165 23783 ne
rect 34165 23780 34428 23783
tri 34428 23780 34436 23788 sw
rect 34165 23775 34436 23780
tri 34165 23770 34170 23775 ne
rect 34170 23772 34436 23775
tri 34436 23772 34444 23780 sw
rect 34170 23770 34444 23772
tri 34170 23762 34178 23770 ne
rect 34178 23764 34444 23770
tri 34444 23764 34452 23772 sw
rect 34178 23762 34452 23764
tri 34178 23754 34186 23762 ne
rect 34186 23756 34452 23762
tri 34452 23756 34460 23764 sw
rect 34186 23754 34460 23756
tri 34186 23746 34194 23754 ne
rect 34194 23748 34460 23754
tri 34460 23748 34468 23756 sw
rect 34194 23746 34468 23748
tri 34194 23738 34202 23746 ne
rect 34202 23740 34468 23746
tri 34468 23740 34476 23748 sw
rect 34202 23738 34476 23740
tri 34202 23730 34210 23738 ne
rect 34210 23732 34476 23738
tri 34476 23732 34484 23740 sw
rect 70802 23732 71000 23790
rect 34210 23730 34484 23732
tri 34210 23722 34218 23730 ne
rect 34218 23724 34484 23730
tri 34484 23724 34492 23732 sw
rect 34218 23722 34492 23724
tri 34218 23714 34226 23722 ne
rect 34226 23716 34492 23722
tri 34492 23716 34500 23724 sw
rect 34226 23714 34500 23716
tri 34226 23706 34234 23714 ne
rect 34234 23708 34500 23714
tri 34500 23708 34508 23716 sw
rect 34234 23706 34508 23708
tri 34234 23698 34242 23706 ne
rect 34242 23704 34508 23706
rect 34242 23698 34374 23704
tri 34242 23690 34250 23698 ne
rect 34250 23690 34374 23698
tri 34250 23682 34258 23690 ne
rect 34258 23682 34374 23690
tri 34258 23674 34266 23682 ne
rect 34266 23674 34374 23682
tri 34266 23666 34274 23674 ne
rect 34274 23666 34374 23674
tri 34274 23658 34282 23666 ne
rect 34282 23658 34374 23666
rect 34420 23700 34508 23704
tri 34508 23700 34516 23708 sw
rect 34420 23692 34516 23700
tri 34516 23692 34524 23700 sw
rect 34420 23684 34524 23692
tri 34524 23684 34532 23692 sw
rect 70802 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23676 34532 23684
tri 34532 23676 34540 23684 sw
rect 34420 23668 34540 23676
tri 34540 23668 34548 23676 sw
rect 34420 23660 34548 23668
tri 34548 23660 34556 23668 sw
rect 34420 23658 34556 23660
tri 34282 23650 34290 23658 ne
rect 34290 23657 34556 23658
tri 34556 23657 34559 23660 sw
rect 34290 23650 34559 23657
tri 34290 23642 34298 23650 ne
rect 34298 23649 34559 23650
tri 34559 23649 34567 23657 sw
rect 34298 23642 34567 23649
tri 34298 23638 34302 23642 ne
rect 34302 23641 34567 23642
tri 34567 23641 34575 23649 sw
rect 34302 23638 34575 23641
tri 34302 23630 34310 23638 ne
rect 34310 23633 34575 23638
tri 34575 23633 34583 23641 sw
rect 34310 23630 34583 23633
tri 34310 23622 34318 23630 ne
rect 34318 23625 34583 23630
tri 34583 23625 34591 23633 sw
rect 70802 23628 71000 23686
rect 34318 23622 34591 23625
tri 34318 23614 34326 23622 ne
rect 34326 23617 34591 23622
tri 34591 23617 34599 23625 sw
rect 34326 23614 34599 23617
tri 34326 23606 34334 23614 ne
rect 34334 23609 34599 23614
tri 34599 23609 34607 23617 sw
rect 34334 23606 34607 23609
tri 34334 23598 34342 23606 ne
rect 34342 23601 34607 23606
tri 34607 23601 34615 23609 sw
rect 34342 23598 34615 23601
tri 34342 23590 34350 23598 ne
rect 34350 23593 34615 23598
tri 34615 23593 34623 23601 sw
rect 34350 23590 34623 23593
tri 34350 23582 34358 23590 ne
rect 34358 23585 34623 23590
tri 34623 23585 34631 23593 sw
rect 34358 23582 34631 23585
tri 34358 23574 34366 23582 ne
rect 34366 23577 34631 23582
tri 34631 23577 34639 23585 sw
rect 70802 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 34366 23574 34639 23577
tri 34366 23571 34369 23574 ne
rect 34369 23572 34639 23574
rect 34369 23571 34506 23572
tri 34369 23563 34377 23571 ne
rect 34377 23563 34506 23571
tri 34377 23555 34385 23563 ne
rect 34385 23555 34506 23563
tri 34385 23547 34393 23555 ne
rect 34393 23547 34506 23555
tri 34393 23539 34401 23547 ne
rect 34401 23539 34506 23547
tri 34401 23531 34409 23539 ne
rect 34409 23531 34506 23539
tri 34409 23523 34417 23531 ne
rect 34417 23526 34506 23531
rect 34552 23571 34639 23572
tri 34639 23571 34645 23577 sw
rect 34552 23563 34645 23571
tri 34645 23563 34653 23571 sw
rect 34552 23555 34653 23563
tri 34653 23555 34661 23563 sw
rect 34552 23547 34661 23555
tri 34661 23547 34669 23555 sw
rect 34552 23539 34669 23547
tri 34669 23539 34677 23547 sw
rect 34552 23531 34677 23539
tri 34677 23531 34685 23539 sw
rect 34552 23526 34685 23531
rect 34417 23523 34685 23526
tri 34685 23523 34693 23531 sw
rect 70802 23524 71000 23582
tri 34417 23515 34425 23523 ne
rect 34425 23515 34693 23523
tri 34693 23515 34701 23523 sw
tri 34425 23507 34433 23515 ne
rect 34433 23507 34701 23515
tri 34701 23507 34709 23515 sw
tri 34433 23499 34441 23507 ne
rect 34441 23499 34709 23507
tri 34709 23499 34717 23507 sw
tri 34441 23491 34449 23499 ne
rect 34449 23491 34717 23499
tri 34717 23491 34725 23499 sw
tri 34449 23483 34457 23491 ne
rect 34457 23483 34725 23491
tri 34725 23483 34733 23491 sw
tri 34457 23475 34465 23483 ne
rect 34465 23475 34733 23483
tri 34733 23475 34741 23483 sw
rect 70802 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
tri 34465 23467 34473 23475 ne
rect 34473 23467 34741 23475
tri 34741 23467 34749 23475 sw
tri 34473 23459 34481 23467 ne
rect 34481 23459 34749 23467
tri 34749 23459 34757 23467 sw
tri 34481 23451 34489 23459 ne
rect 34489 23451 34757 23459
tri 34757 23451 34765 23459 sw
tri 34489 23443 34497 23451 ne
rect 34497 23443 34765 23451
tri 34765 23443 34773 23451 sw
tri 34497 23435 34505 23443 ne
rect 34505 23440 34773 23443
rect 34505 23435 34638 23440
tri 34505 23433 34507 23435 ne
rect 34507 23433 34638 23435
tri 34507 23425 34515 23433 ne
rect 34515 23425 34638 23433
tri 34515 23417 34523 23425 ne
rect 34523 23417 34638 23425
tri 34523 23409 34531 23417 ne
rect 34531 23409 34638 23417
tri 34531 23401 34539 23409 ne
rect 34539 23401 34638 23409
tri 34539 23393 34547 23401 ne
rect 34547 23394 34638 23401
rect 34684 23435 34773 23440
tri 34773 23435 34781 23443 sw
rect 34684 23433 34781 23435
tri 34781 23433 34783 23435 sw
rect 34684 23425 34783 23433
tri 34783 23425 34791 23433 sw
rect 34684 23417 34791 23425
tri 34791 23417 34799 23425 sw
rect 70802 23420 71000 23478
rect 34684 23409 34799 23417
tri 34799 23409 34807 23417 sw
rect 34684 23401 34807 23409
tri 34807 23401 34815 23409 sw
rect 34684 23394 34815 23401
rect 34547 23393 34815 23394
tri 34815 23393 34823 23401 sw
tri 34547 23385 34555 23393 ne
rect 34555 23385 34823 23393
tri 34823 23385 34831 23393 sw
tri 34555 23377 34563 23385 ne
rect 34563 23377 34831 23385
tri 34831 23377 34839 23385 sw
tri 34563 23369 34571 23377 ne
rect 34571 23369 34839 23377
tri 34839 23369 34847 23377 sw
rect 70802 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34571 23361 34579 23369 ne
rect 34579 23361 34847 23369
tri 34847 23361 34855 23369 sw
tri 34579 23353 34587 23361 ne
rect 34587 23353 34855 23361
tri 34855 23353 34863 23361 sw
tri 34587 23345 34595 23353 ne
rect 34595 23345 34863 23353
tri 34863 23345 34871 23353 sw
tri 34595 23337 34603 23345 ne
rect 34603 23337 34871 23345
tri 34871 23337 34879 23345 sw
tri 34603 23329 34611 23337 ne
rect 34611 23329 34879 23337
tri 34879 23329 34887 23337 sw
tri 34611 23321 34619 23329 ne
rect 34619 23321 34887 23329
tri 34887 23321 34895 23329 sw
tri 34619 23313 34627 23321 ne
rect 34627 23313 34895 23321
tri 34895 23313 34903 23321 sw
rect 70802 23316 71000 23374
tri 34627 23309 34631 23313 ne
rect 34631 23309 34903 23313
tri 34903 23309 34907 23313 sw
tri 34631 23305 34635 23309 ne
rect 34635 23308 34907 23309
rect 34635 23305 34770 23308
tri 34635 23297 34643 23305 ne
rect 34643 23297 34770 23305
tri 34643 23289 34651 23297 ne
rect 34651 23289 34770 23297
tri 34651 23281 34659 23289 ne
rect 34659 23281 34770 23289
tri 34659 23273 34667 23281 ne
rect 34667 23273 34770 23281
tri 34667 23265 34675 23273 ne
rect 34675 23265 34770 23273
tri 34675 23257 34683 23265 ne
rect 34683 23262 34770 23265
rect 34816 23305 34907 23308
tri 34907 23305 34911 23309 sw
rect 34816 23297 34911 23305
tri 34911 23297 34919 23305 sw
rect 34816 23289 34919 23297
tri 34919 23289 34927 23297 sw
rect 34816 23281 34927 23289
tri 34927 23281 34935 23289 sw
rect 34816 23273 34935 23281
tri 34935 23273 34943 23281 sw
rect 34816 23265 34943 23273
tri 34943 23265 34951 23273 sw
rect 70802 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 34816 23262 34951 23265
rect 34683 23257 34951 23262
tri 34951 23257 34959 23265 sw
tri 34683 23249 34691 23257 ne
rect 34691 23249 34959 23257
tri 34959 23249 34967 23257 sw
tri 34691 23241 34699 23249 ne
rect 34699 23241 34967 23249
tri 34967 23241 34975 23249 sw
tri 34699 23233 34707 23241 ne
rect 34707 23233 34975 23241
tri 34975 23233 34983 23241 sw
tri 34707 23225 34715 23233 ne
rect 34715 23225 34983 23233
tri 34983 23225 34991 23233 sw
tri 34715 23217 34723 23225 ne
rect 34723 23217 34991 23225
tri 34991 23217 34999 23225 sw
tri 34723 23209 34731 23217 ne
rect 34731 23209 34999 23217
tri 34999 23209 35007 23217 sw
rect 70802 23212 71000 23270
tri 34731 23201 34739 23209 ne
rect 34739 23201 35007 23209
tri 35007 23201 35015 23209 sw
tri 34739 23193 34747 23201 ne
rect 34747 23193 35015 23201
tri 35015 23193 35023 23201 sw
tri 34747 23185 34755 23193 ne
rect 34755 23190 35023 23193
tri 35023 23190 35026 23193 sw
rect 34755 23185 35026 23190
tri 34755 23177 34763 23185 ne
rect 34763 23182 35026 23185
tri 35026 23182 35034 23190 sw
rect 34763 23177 35034 23182
tri 34763 23169 34771 23177 ne
rect 34771 23176 35034 23177
rect 34771 23169 34902 23176
tri 34771 23166 34774 23169 ne
rect 34774 23166 34902 23169
tri 34774 23158 34782 23166 ne
rect 34782 23158 34902 23166
tri 34782 23150 34790 23158 ne
rect 34790 23150 34902 23158
tri 34790 23142 34798 23150 ne
rect 34798 23142 34902 23150
tri 34798 23134 34806 23142 ne
rect 34806 23134 34902 23142
tri 34806 23126 34814 23134 ne
rect 34814 23130 34902 23134
rect 34948 23174 35034 23176
tri 35034 23174 35042 23182 sw
rect 34948 23166 35042 23174
tri 35042 23166 35050 23174 sw
rect 70802 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 34948 23158 35050 23166
tri 35050 23158 35058 23166 sw
rect 34948 23150 35058 23158
tri 35058 23150 35066 23158 sw
rect 34948 23142 35066 23150
tri 35066 23142 35074 23150 sw
rect 34948 23134 35074 23142
tri 35074 23134 35082 23142 sw
rect 34948 23130 35082 23134
rect 34814 23126 35082 23130
tri 35082 23126 35090 23134 sw
tri 34814 23118 34822 23126 ne
rect 34822 23118 35090 23126
tri 35090 23118 35098 23126 sw
tri 34822 23110 34830 23118 ne
rect 34830 23110 35098 23118
tri 35098 23110 35106 23118 sw
tri 34830 23102 34838 23110 ne
rect 34838 23102 35106 23110
tri 35106 23102 35114 23110 sw
rect 70802 23108 71000 23166
tri 34838 23094 34846 23102 ne
rect 34846 23094 35114 23102
tri 35114 23094 35122 23102 sw
tri 34846 23086 34854 23094 ne
rect 34854 23086 35122 23094
tri 35122 23086 35130 23094 sw
tri 34854 23078 34862 23086 ne
rect 34862 23078 35130 23086
tri 35130 23078 35138 23086 sw
tri 34862 23070 34870 23078 ne
rect 34870 23070 35138 23078
tri 35138 23070 35146 23078 sw
tri 34870 23062 34878 23070 ne
rect 34878 23062 35146 23070
tri 35146 23062 35154 23070 sw
rect 70802 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
tri 34878 23054 34886 23062 ne
rect 34886 23054 35154 23062
tri 35154 23054 35162 23062 sw
tri 34886 23046 34894 23054 ne
rect 34894 23047 35162 23054
tri 35162 23047 35169 23054 sw
rect 34894 23046 35169 23047
tri 34894 23038 34902 23046 ne
rect 34902 23044 35169 23046
rect 34902 23038 35034 23044
tri 34902 23031 34909 23038 ne
rect 34909 23031 35034 23038
tri 34909 23029 34911 23031 ne
rect 34911 23029 35034 23031
tri 34911 23023 34917 23029 ne
rect 34917 23023 35034 23029
tri 34917 23015 34925 23023 ne
rect 34925 23015 35034 23023
tri 34925 23007 34933 23015 ne
rect 34933 23007 35034 23015
tri 34933 22999 34941 23007 ne
rect 34941 22999 35034 23007
tri 34941 22991 34949 22999 ne
rect 34949 22998 35034 22999
rect 35080 23039 35169 23044
tri 35169 23039 35177 23047 sw
rect 35080 23031 35177 23039
tri 35177 23031 35185 23039 sw
rect 35080 23023 35185 23031
tri 35185 23023 35193 23031 sw
rect 35080 23015 35193 23023
tri 35193 23015 35201 23023 sw
rect 35080 23007 35201 23015
tri 35201 23007 35209 23015 sw
rect 35080 22999 35209 23007
tri 35209 22999 35217 23007 sw
rect 70802 23004 71000 23062
rect 35080 22998 35217 22999
rect 34949 22991 35217 22998
tri 35217 22991 35225 22999 sw
tri 34949 22983 34957 22991 ne
rect 34957 22983 35225 22991
tri 35225 22983 35233 22991 sw
tri 34957 22979 34961 22983 ne
rect 34961 22979 35233 22983
tri 35233 22979 35237 22983 sw
tri 34961 22971 34969 22979 ne
rect 34969 22971 35237 22979
tri 35237 22971 35245 22979 sw
tri 34969 22963 34977 22971 ne
rect 34977 22963 35245 22971
tri 35245 22963 35253 22971 sw
tri 34977 22955 34985 22963 ne
rect 34985 22955 35253 22963
tri 35253 22955 35261 22963 sw
rect 70802 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 34985 22947 34993 22955 ne
rect 34993 22947 35261 22955
tri 35261 22947 35269 22955 sw
tri 34993 22939 35001 22947 ne
rect 35001 22939 35269 22947
tri 35269 22939 35277 22947 sw
tri 35001 22931 35009 22939 ne
rect 35009 22931 35277 22939
tri 35277 22931 35285 22939 sw
tri 35009 22923 35017 22931 ne
rect 35017 22923 35285 22931
tri 35285 22923 35293 22931 sw
tri 35017 22915 35025 22923 ne
rect 35025 22915 35293 22923
tri 35293 22915 35301 22923 sw
tri 35025 22907 35033 22915 ne
rect 35033 22912 35301 22915
rect 35033 22907 35166 22912
tri 35033 22899 35041 22907 ne
rect 35041 22899 35166 22907
tri 35041 22891 35049 22899 ne
rect 35049 22891 35166 22899
tri 35049 22883 35057 22891 ne
rect 35057 22883 35166 22891
tri 35057 22875 35065 22883 ne
rect 35065 22875 35166 22883
tri 35065 22867 35073 22875 ne
rect 35073 22867 35166 22875
tri 35073 22859 35081 22867 ne
rect 35081 22866 35166 22867
rect 35212 22907 35301 22912
tri 35301 22907 35309 22915 sw
rect 35212 22899 35309 22907
tri 35309 22899 35317 22907 sw
rect 70802 22900 71000 22958
rect 35212 22891 35317 22899
tri 35317 22891 35325 22899 sw
rect 35212 22883 35325 22891
tri 35325 22883 35333 22891 sw
rect 35212 22875 35333 22883
tri 35333 22875 35341 22883 sw
rect 35212 22874 35341 22875
tri 35341 22874 35342 22875 sw
rect 35212 22866 35342 22874
tri 35342 22866 35350 22874 sw
rect 35081 22859 35350 22866
tri 35081 22854 35086 22859 ne
rect 35086 22858 35350 22859
tri 35350 22858 35358 22866 sw
rect 35086 22854 35358 22858
tri 35086 22846 35094 22854 ne
rect 35094 22850 35358 22854
tri 35358 22850 35366 22858 sw
rect 70802 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
rect 35094 22846 35366 22850
tri 35094 22838 35102 22846 ne
rect 35102 22842 35366 22846
tri 35366 22842 35374 22850 sw
rect 35102 22838 35374 22842
tri 35102 22830 35110 22838 ne
rect 35110 22834 35374 22838
tri 35374 22834 35382 22842 sw
rect 35110 22830 35382 22834
tri 35110 22822 35118 22830 ne
rect 35118 22826 35382 22830
tri 35382 22826 35390 22834 sw
rect 35118 22822 35390 22826
tri 35118 22814 35126 22822 ne
rect 35126 22818 35390 22822
tri 35390 22818 35398 22826 sw
rect 35126 22814 35398 22818
tri 35126 22806 35134 22814 ne
rect 35134 22810 35398 22814
tri 35398 22810 35406 22818 sw
rect 35134 22806 35406 22810
tri 35134 22798 35142 22806 ne
rect 35142 22802 35406 22806
tri 35406 22802 35414 22810 sw
rect 35142 22798 35414 22802
tri 35142 22790 35150 22798 ne
rect 35150 22794 35414 22798
tri 35414 22794 35422 22802 sw
rect 70802 22796 71000 22854
rect 35150 22790 35422 22794
tri 35150 22782 35158 22790 ne
rect 35158 22786 35422 22790
tri 35422 22786 35430 22794 sw
rect 35158 22782 35430 22786
tri 35158 22774 35166 22782 ne
rect 35166 22780 35430 22782
rect 35166 22774 35298 22780
tri 35166 22766 35174 22774 ne
rect 35174 22766 35298 22774
tri 35174 22758 35182 22766 ne
rect 35182 22758 35298 22766
tri 35182 22755 35185 22758 ne
rect 35185 22755 35298 22758
tri 35185 22747 35193 22755 ne
rect 35193 22747 35298 22755
tri 35193 22739 35201 22747 ne
rect 35201 22739 35298 22747
tri 35201 22731 35209 22739 ne
rect 35209 22734 35298 22739
rect 35344 22778 35430 22780
tri 35430 22778 35438 22786 sw
rect 35344 22770 35438 22778
tri 35438 22770 35446 22778 sw
rect 35344 22763 35446 22770
tri 35446 22763 35453 22770 sw
rect 35344 22755 35453 22763
tri 35453 22755 35461 22763 sw
rect 35344 22747 35461 22755
tri 35461 22747 35469 22755 sw
rect 70802 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 35344 22739 35469 22747
tri 35469 22739 35477 22747 sw
rect 35344 22734 35477 22739
rect 35209 22731 35477 22734
tri 35477 22731 35485 22739 sw
tri 35209 22723 35217 22731 ne
rect 35217 22723 35485 22731
tri 35485 22723 35493 22731 sw
tri 35217 22715 35225 22723 ne
rect 35225 22715 35493 22723
tri 35493 22715 35501 22723 sw
tri 35225 22707 35233 22715 ne
rect 35233 22707 35501 22715
tri 35501 22707 35509 22715 sw
tri 35233 22699 35241 22707 ne
rect 35241 22699 35509 22707
tri 35509 22699 35517 22707 sw
tri 35241 22691 35249 22699 ne
rect 35249 22695 35517 22699
tri 35517 22695 35521 22699 sw
rect 35249 22691 35521 22695
tri 35249 22683 35257 22691 ne
rect 35257 22687 35521 22691
tri 35521 22687 35529 22695 sw
rect 70802 22692 71000 22750
rect 35257 22683 35529 22687
tri 35257 22675 35265 22683 ne
rect 35265 22679 35529 22683
tri 35529 22679 35537 22687 sw
rect 35265 22675 35537 22679
tri 35265 22667 35273 22675 ne
rect 35273 22671 35537 22675
tri 35537 22671 35545 22679 sw
rect 35273 22667 35545 22671
tri 35273 22659 35281 22667 ne
rect 35281 22663 35545 22667
tri 35545 22663 35553 22671 sw
rect 35281 22659 35553 22663
tri 35281 22651 35289 22659 ne
rect 35289 22655 35553 22659
tri 35553 22655 35561 22663 sw
rect 35289 22651 35561 22655
tri 35289 22643 35297 22651 ne
rect 35297 22648 35561 22651
rect 35297 22643 35430 22648
tri 35297 22635 35305 22643 ne
rect 35305 22635 35430 22643
tri 35305 22627 35313 22635 ne
rect 35313 22627 35430 22635
tri 35313 22619 35321 22627 ne
rect 35321 22619 35430 22627
tri 35321 22611 35329 22619 ne
rect 35329 22611 35430 22619
tri 35329 22603 35337 22611 ne
rect 35337 22603 35430 22611
tri 35337 22595 35345 22603 ne
rect 35345 22602 35430 22603
rect 35476 22647 35561 22648
tri 35561 22647 35569 22655 sw
rect 35476 22639 35569 22647
tri 35569 22639 35577 22647 sw
rect 70802 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22631 35577 22639
tri 35577 22631 35585 22639 sw
rect 35476 22623 35585 22631
tri 35585 22623 35593 22631 sw
rect 35476 22615 35593 22623
tri 35593 22615 35601 22623 sw
rect 35476 22607 35601 22615
tri 35601 22607 35609 22615 sw
rect 35476 22602 35609 22607
rect 35345 22599 35609 22602
tri 35609 22599 35617 22607 sw
rect 35345 22598 35617 22599
tri 35617 22598 35618 22599 sw
rect 35345 22595 35618 22598
tri 35345 22587 35353 22595 ne
rect 35353 22590 35618 22595
tri 35618 22590 35626 22598 sw
rect 35353 22587 35626 22590
tri 35353 22582 35358 22587 ne
rect 35358 22582 35626 22587
tri 35626 22582 35634 22590 sw
rect 70802 22588 71000 22646
tri 35358 22574 35366 22582 ne
rect 35366 22574 35634 22582
tri 35634 22574 35642 22582 sw
tri 35366 22566 35374 22574 ne
rect 35374 22566 35642 22574
tri 35642 22566 35650 22574 sw
tri 35374 22558 35382 22566 ne
rect 35382 22558 35650 22566
tri 35650 22558 35658 22566 sw
tri 35382 22550 35390 22558 ne
rect 35390 22550 35658 22558
tri 35658 22550 35666 22558 sw
tri 35390 22542 35398 22550 ne
rect 35398 22542 35666 22550
tri 35666 22542 35674 22550 sw
rect 70802 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35398 22534 35406 22542 ne
rect 35406 22534 35674 22542
tri 35674 22534 35682 22542 sw
tri 35406 22526 35414 22534 ne
rect 35414 22526 35682 22534
tri 35682 22526 35690 22534 sw
tri 35414 22518 35422 22526 ne
rect 35422 22518 35690 22526
tri 35690 22518 35698 22526 sw
tri 35422 22510 35430 22518 ne
rect 35430 22516 35698 22518
rect 35430 22510 35562 22516
tri 35430 22502 35438 22510 ne
rect 35438 22502 35562 22510
tri 35438 22494 35446 22502 ne
rect 35446 22494 35562 22502
tri 35446 22486 35454 22494 ne
rect 35454 22486 35562 22494
tri 35454 22483 35457 22486 ne
rect 35457 22483 35562 22486
tri 35457 22475 35465 22483 ne
rect 35465 22475 35562 22483
tri 35465 22467 35473 22475 ne
rect 35473 22470 35562 22475
rect 35608 22511 35698 22516
tri 35698 22511 35705 22518 sw
rect 35608 22503 35705 22511
tri 35705 22503 35713 22511 sw
rect 35608 22495 35713 22503
tri 35713 22495 35721 22503 sw
rect 35608 22487 35721 22495
tri 35721 22487 35729 22495 sw
rect 35608 22479 35729 22487
tri 35729 22479 35737 22487 sw
rect 70802 22484 71000 22542
rect 35608 22475 35737 22479
tri 35737 22475 35741 22479 sw
rect 35608 22470 35741 22475
rect 35473 22467 35741 22470
tri 35741 22467 35749 22475 sw
tri 35473 22459 35481 22467 ne
rect 35481 22459 35749 22467
tri 35749 22459 35757 22467 sw
tri 35481 22451 35489 22459 ne
rect 35489 22451 35757 22459
tri 35757 22451 35765 22459 sw
tri 35489 22443 35497 22451 ne
rect 35497 22443 35765 22451
tri 35765 22443 35773 22451 sw
tri 35497 22435 35505 22443 ne
rect 35505 22435 35773 22443
tri 35773 22435 35781 22443 sw
rect 70802 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35505 22427 35513 22435 ne
rect 35513 22427 35781 22435
tri 35781 22427 35789 22435 sw
tri 35513 22419 35521 22427 ne
rect 35521 22423 35789 22427
tri 35789 22423 35793 22427 sw
rect 35521 22419 35793 22423
tri 35521 22415 35525 22419 ne
rect 35525 22415 35793 22419
tri 35793 22415 35801 22423 sw
tri 35525 22407 35533 22415 ne
rect 35533 22407 35801 22415
tri 35801 22407 35809 22415 sw
tri 35533 22399 35541 22407 ne
rect 35541 22399 35809 22407
tri 35809 22399 35817 22407 sw
tri 35541 22391 35549 22399 ne
rect 35549 22391 35817 22399
tri 35817 22391 35825 22399 sw
tri 35549 22383 35557 22391 ne
rect 35557 22384 35825 22391
rect 35557 22383 35694 22384
tri 35557 22375 35565 22383 ne
rect 35565 22375 35694 22383
tri 35565 22367 35573 22375 ne
rect 35573 22367 35694 22375
tri 35573 22359 35581 22367 ne
rect 35581 22359 35694 22367
tri 35581 22351 35589 22359 ne
rect 35589 22351 35694 22359
tri 35589 22343 35597 22351 ne
rect 35597 22343 35694 22351
tri 35597 22335 35605 22343 ne
rect 35605 22338 35694 22343
rect 35740 22383 35825 22384
tri 35825 22383 35833 22391 sw
rect 35740 22375 35833 22383
tri 35833 22375 35841 22383 sw
rect 70802 22380 71000 22438
rect 35740 22367 35841 22375
tri 35841 22367 35849 22375 sw
rect 35740 22359 35849 22367
tri 35849 22359 35857 22367 sw
rect 35740 22351 35857 22359
tri 35857 22351 35865 22359 sw
rect 35740 22343 35865 22351
tri 35865 22343 35873 22351 sw
rect 35740 22338 35873 22343
rect 35605 22335 35873 22338
tri 35873 22335 35881 22343 sw
tri 35605 22327 35613 22335 ne
rect 35613 22327 35881 22335
tri 35881 22327 35889 22335 sw
rect 70802 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35613 22319 35621 22327 ne
rect 35621 22319 35889 22327
tri 35889 22319 35897 22327 sw
tri 35621 22311 35629 22319 ne
rect 35629 22311 35897 22319
tri 35897 22311 35905 22319 sw
tri 35629 22303 35637 22311 ne
rect 35637 22303 35905 22311
tri 35905 22303 35913 22311 sw
tri 35637 22299 35641 22303 ne
rect 35641 22299 35913 22303
tri 35913 22299 35917 22303 sw
tri 35641 22291 35649 22299 ne
rect 35649 22291 35917 22299
tri 35917 22291 35925 22299 sw
tri 35649 22283 35657 22291 ne
rect 35657 22283 35925 22291
tri 35925 22283 35933 22291 sw
tri 35657 22275 35665 22283 ne
rect 35665 22275 35933 22283
tri 35933 22275 35941 22283 sw
rect 70802 22276 71000 22334
tri 35665 22267 35673 22275 ne
rect 35673 22267 35941 22275
tri 35941 22267 35949 22275 sw
tri 35673 22259 35681 22267 ne
rect 35681 22259 35949 22267
tri 35949 22259 35957 22267 sw
tri 35681 22251 35689 22259 ne
rect 35689 22252 35957 22259
rect 35689 22251 35826 22252
tri 35689 22243 35697 22251 ne
rect 35697 22243 35826 22251
tri 35697 22235 35705 22243 ne
rect 35705 22235 35826 22243
tri 35705 22227 35713 22235 ne
rect 35713 22227 35826 22235
tri 35713 22219 35721 22227 ne
rect 35721 22219 35826 22227
tri 35721 22211 35729 22219 ne
rect 35729 22211 35826 22219
tri 35729 22203 35737 22211 ne
rect 35737 22206 35826 22211
rect 35872 22251 35957 22252
tri 35957 22251 35965 22259 sw
rect 35872 22243 35965 22251
tri 35965 22243 35973 22251 sw
rect 35872 22235 35973 22243
tri 35973 22235 35981 22243 sw
rect 35872 22227 35981 22235
tri 35981 22227 35989 22235 sw
rect 70802 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22219 35989 22227
tri 35989 22219 35997 22227 sw
rect 35872 22211 35997 22219
tri 35997 22211 36005 22219 sw
rect 35872 22206 36005 22211
rect 35737 22203 36005 22206
tri 36005 22203 36013 22211 sw
tri 35737 22195 35745 22203 ne
rect 35745 22195 36013 22203
tri 36013 22195 36021 22203 sw
tri 35745 22187 35753 22195 ne
rect 35753 22187 36021 22195
tri 36021 22187 36029 22195 sw
tri 35753 22179 35761 22187 ne
rect 35761 22179 36029 22187
tri 36029 22179 36037 22187 sw
tri 35761 22171 35769 22179 ne
rect 35769 22171 36037 22179
tri 36037 22171 36045 22179 sw
rect 70802 22172 71000 22230
tri 35769 22163 35777 22171 ne
rect 35777 22165 36045 22171
tri 36045 22165 36051 22171 sw
rect 35777 22163 36051 22165
tri 35777 22155 35785 22163 ne
rect 35785 22157 36051 22163
tri 36051 22157 36059 22165 sw
rect 35785 22155 36059 22157
tri 35785 22147 35793 22155 ne
rect 35793 22149 36059 22155
tri 36059 22149 36067 22157 sw
rect 35793 22147 36067 22149
tri 35793 22139 35801 22147 ne
rect 35801 22141 36067 22147
tri 36067 22141 36075 22149 sw
rect 35801 22139 36075 22141
tri 35801 22131 35809 22139 ne
rect 35809 22133 36075 22139
tri 36075 22133 36083 22141 sw
rect 35809 22131 36083 22133
tri 35809 22123 35817 22131 ne
rect 35817 22125 36083 22131
tri 36083 22125 36091 22133 sw
rect 70802 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 35817 22123 36091 22125
tri 35817 22115 35825 22123 ne
rect 35825 22120 36091 22123
rect 35825 22115 35958 22120
tri 35825 22107 35833 22115 ne
rect 35833 22107 35958 22115
tri 35833 22099 35841 22107 ne
rect 35841 22099 35958 22107
tri 35841 22091 35849 22099 ne
rect 35849 22091 35958 22099
tri 35849 22083 35857 22091 ne
rect 35857 22083 35958 22091
tri 35857 22075 35865 22083 ne
rect 35865 22075 35958 22083
tri 35865 22067 35873 22075 ne
rect 35873 22074 35958 22075
rect 36004 22117 36091 22120
tri 36091 22117 36099 22125 sw
rect 36004 22109 36099 22117
tri 36099 22109 36107 22117 sw
rect 36004 22101 36107 22109
tri 36107 22101 36115 22109 sw
rect 36004 22093 36115 22101
tri 36115 22093 36123 22101 sw
rect 36004 22085 36123 22093
tri 36123 22085 36131 22093 sw
rect 36004 22077 36131 22085
tri 36131 22077 36139 22085 sw
rect 36004 22074 36139 22077
rect 35873 22069 36139 22074
tri 36139 22069 36147 22077 sw
rect 35873 22067 36147 22069
tri 35873 22059 35881 22067 ne
rect 35881 22061 36147 22067
tri 36147 22061 36155 22069 sw
rect 70802 22068 71000 22126
rect 35881 22059 36155 22061
tri 35881 22051 35889 22059 ne
rect 35889 22055 36155 22059
tri 36155 22055 36161 22061 sw
rect 35889 22051 36161 22055
tri 35889 22050 35890 22051 ne
rect 35890 22050 36161 22051
tri 35890 22042 35898 22050 ne
rect 35898 22047 36161 22050
tri 36161 22047 36169 22055 sw
rect 35898 22042 36169 22047
tri 35898 22034 35906 22042 ne
rect 35906 22039 36169 22042
tri 36169 22039 36177 22047 sw
rect 35906 22034 36177 22039
tri 35906 22026 35914 22034 ne
rect 35914 22031 36177 22034
tri 36177 22031 36185 22039 sw
rect 35914 22026 36185 22031
tri 35914 22018 35922 22026 ne
rect 35922 22023 36185 22026
tri 36185 22023 36193 22031 sw
rect 35922 22018 36193 22023
tri 35922 22010 35930 22018 ne
rect 35930 22015 36193 22018
tri 36193 22015 36201 22023 sw
rect 70802 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
rect 35930 22010 36201 22015
tri 35930 22002 35938 22010 ne
rect 35938 22007 36201 22010
tri 36201 22007 36209 22015 sw
rect 35938 22002 36209 22007
tri 35938 21994 35946 22002 ne
rect 35946 21999 36209 22002
tri 36209 21999 36217 22007 sw
rect 35946 21994 36217 21999
tri 35946 21986 35954 21994 ne
rect 35954 21991 36217 21994
tri 36217 21991 36225 21999 sw
rect 35954 21988 36225 21991
rect 35954 21986 36090 21988
tri 35954 21978 35962 21986 ne
rect 35962 21978 36090 21986
tri 35962 21970 35970 21978 ne
rect 35970 21970 36090 21978
tri 35970 21962 35978 21970 ne
rect 35978 21962 36090 21970
tri 35978 21954 35986 21962 ne
rect 35986 21954 36090 21962
tri 35986 21946 35994 21954 ne
rect 35994 21946 36090 21954
tri 35994 21938 36002 21946 ne
rect 36002 21942 36090 21946
rect 36136 21983 36225 21988
tri 36225 21983 36233 21991 sw
rect 36136 21978 36233 21983
tri 36233 21978 36238 21983 sw
rect 36136 21975 36238 21978
tri 36238 21975 36241 21978 sw
rect 36136 21967 36241 21975
tri 36241 21967 36249 21975 sw
rect 36136 21959 36249 21967
tri 36249 21959 36257 21967 sw
rect 70802 21964 71000 22022
rect 36136 21951 36257 21959
tri 36257 21951 36265 21959 sw
rect 36136 21943 36265 21951
tri 36265 21943 36273 21951 sw
rect 36136 21942 36273 21943
rect 36002 21938 36273 21942
tri 36002 21930 36010 21938 ne
rect 36010 21935 36273 21938
tri 36273 21935 36281 21943 sw
rect 36010 21934 36281 21935
tri 36281 21934 36282 21935 sw
rect 36010 21930 36282 21934
tri 36010 21924 36016 21930 ne
rect 36016 21926 36282 21930
tri 36282 21926 36290 21934 sw
rect 36016 21924 36290 21926
tri 36016 21916 36024 21924 ne
rect 36024 21918 36290 21924
tri 36290 21918 36298 21926 sw
rect 70802 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36024 21916 36298 21918
tri 36024 21908 36032 21916 ne
rect 36032 21910 36298 21916
tri 36298 21910 36306 21918 sw
rect 36032 21908 36306 21910
tri 36032 21900 36040 21908 ne
rect 36040 21902 36306 21908
tri 36306 21902 36314 21910 sw
rect 36040 21900 36314 21902
tri 36040 21892 36048 21900 ne
rect 36048 21894 36314 21900
tri 36314 21894 36322 21902 sw
rect 36048 21892 36322 21894
tri 36048 21884 36056 21892 ne
rect 36056 21886 36322 21892
tri 36322 21886 36330 21894 sw
rect 36056 21884 36330 21886
tri 36056 21876 36064 21884 ne
rect 36064 21878 36330 21884
tri 36330 21878 36338 21886 sw
rect 36064 21876 36338 21878
tri 36064 21868 36072 21876 ne
rect 36072 21870 36338 21876
tri 36338 21870 36346 21878 sw
rect 36072 21868 36346 21870
tri 36072 21860 36080 21868 ne
rect 36080 21862 36346 21868
tri 36346 21862 36354 21870 sw
rect 36080 21860 36354 21862
tri 36080 21852 36088 21860 ne
rect 36088 21856 36354 21860
rect 36088 21852 36222 21856
tri 36088 21844 36096 21852 ne
rect 36096 21844 36222 21852
tri 36096 21836 36104 21844 ne
rect 36104 21836 36222 21844
tri 36104 21828 36112 21836 ne
rect 36112 21828 36222 21836
tri 36112 21820 36120 21828 ne
rect 36120 21820 36222 21828
tri 36120 21812 36128 21820 ne
rect 36128 21812 36222 21820
tri 36128 21804 36136 21812 ne
rect 36136 21810 36222 21812
rect 36268 21854 36354 21856
tri 36354 21854 36362 21862 sw
rect 70802 21860 71000 21918
rect 36268 21846 36362 21854
tri 36362 21846 36370 21854 sw
rect 36268 21838 36370 21846
tri 36370 21838 36378 21846 sw
rect 36268 21830 36378 21838
tri 36378 21830 36386 21838 sw
rect 36268 21822 36386 21830
tri 36386 21822 36394 21830 sw
rect 36268 21815 36394 21822
tri 36394 21815 36401 21822 sw
rect 36268 21810 36401 21815
rect 36136 21807 36401 21810
tri 36401 21807 36409 21815 sw
rect 70802 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 36136 21804 36409 21807
tri 36136 21798 36142 21804 ne
rect 36142 21799 36409 21804
tri 36409 21799 36417 21807 sw
rect 36142 21798 36417 21799
tri 36142 21790 36150 21798 ne
rect 36150 21791 36417 21798
tri 36417 21791 36425 21799 sw
rect 36150 21790 36425 21791
tri 36150 21782 36158 21790 ne
rect 36158 21783 36425 21790
tri 36425 21783 36433 21791 sw
rect 36158 21782 36433 21783
tri 36158 21774 36166 21782 ne
rect 36166 21775 36433 21782
tri 36433 21775 36441 21783 sw
rect 36166 21774 36441 21775
tri 36166 21766 36174 21774 ne
rect 36174 21767 36441 21774
tri 36441 21767 36449 21775 sw
rect 36174 21766 36449 21767
tri 36174 21758 36182 21766 ne
rect 36182 21759 36449 21766
tri 36449 21759 36457 21767 sw
rect 36182 21758 36457 21759
tri 36182 21750 36190 21758 ne
rect 36190 21751 36457 21758
tri 36457 21751 36465 21759 sw
rect 70802 21756 71000 21814
rect 36190 21750 36465 21751
tri 36190 21742 36198 21750 ne
rect 36198 21743 36465 21750
tri 36465 21743 36473 21751 sw
rect 36198 21742 36473 21743
tri 36198 21734 36206 21742 ne
rect 36206 21735 36473 21742
tri 36473 21735 36481 21743 sw
rect 36206 21734 36481 21735
tri 36206 21726 36214 21734 ne
rect 36214 21727 36481 21734
tri 36481 21727 36489 21735 sw
rect 36214 21726 36489 21727
tri 36214 21718 36222 21726 ne
rect 36222 21724 36489 21726
rect 36222 21718 36354 21724
tri 36222 21710 36230 21718 ne
rect 36230 21710 36354 21718
tri 36230 21707 36233 21710 ne
rect 36233 21707 36354 21710
tri 36233 21699 36241 21707 ne
rect 36241 21699 36354 21707
tri 36241 21691 36249 21699 ne
rect 36249 21691 36354 21699
tri 36249 21683 36257 21691 ne
rect 36257 21683 36354 21691
tri 36257 21675 36265 21683 ne
rect 36265 21678 36354 21683
rect 36400 21719 36489 21724
tri 36489 21719 36497 21727 sw
rect 36400 21715 36497 21719
tri 36497 21715 36501 21719 sw
rect 36400 21707 36501 21715
tri 36501 21707 36509 21715 sw
rect 70802 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 36400 21699 36509 21707
tri 36509 21699 36517 21707 sw
rect 36400 21691 36517 21699
tri 36517 21691 36525 21699 sw
rect 36400 21683 36525 21691
tri 36525 21683 36533 21691 sw
rect 36400 21678 36533 21683
rect 36265 21675 36533 21678
tri 36533 21675 36541 21683 sw
tri 36265 21667 36273 21675 ne
rect 36273 21667 36541 21675
tri 36541 21667 36549 21675 sw
tri 36273 21659 36281 21667 ne
rect 36281 21659 36549 21667
tri 36549 21659 36557 21667 sw
tri 36281 21651 36289 21659 ne
rect 36289 21651 36557 21659
tri 36557 21651 36565 21659 sw
rect 70802 21652 71000 21710
tri 36289 21648 36292 21651 ne
rect 36292 21648 36565 21651
tri 36565 21648 36568 21651 sw
tri 36292 21640 36300 21648 ne
rect 36300 21640 36568 21648
tri 36568 21640 36576 21648 sw
tri 36300 21632 36308 21640 ne
rect 36308 21632 36576 21640
tri 36576 21632 36584 21640 sw
tri 36308 21624 36316 21632 ne
rect 36316 21624 36584 21632
tri 36584 21624 36592 21632 sw
tri 36316 21616 36324 21624 ne
rect 36324 21616 36592 21624
tri 36592 21616 36600 21624 sw
tri 36324 21608 36332 21616 ne
rect 36332 21608 36600 21616
tri 36600 21608 36608 21616 sw
tri 36332 21600 36340 21608 ne
rect 36340 21600 36608 21608
tri 36608 21600 36616 21608 sw
rect 70802 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
tri 36340 21592 36348 21600 ne
rect 36348 21592 36616 21600
tri 36616 21592 36624 21600 sw
tri 36348 21584 36356 21592 ne
rect 36356 21584 36486 21592
tri 36356 21576 36364 21584 ne
rect 36364 21576 36486 21584
tri 36364 21568 36372 21576 ne
rect 36372 21568 36486 21576
tri 36372 21560 36380 21568 ne
rect 36380 21560 36486 21568
tri 36380 21552 36388 21560 ne
rect 36388 21552 36486 21560
tri 36388 21544 36396 21552 ne
rect 36396 21546 36486 21552
rect 36532 21584 36624 21592
tri 36624 21584 36632 21592 sw
rect 36532 21576 36632 21584
tri 36632 21576 36640 21584 sw
rect 36532 21568 36640 21576
tri 36640 21568 36648 21576 sw
rect 36532 21560 36648 21568
tri 36648 21560 36656 21568 sw
rect 36532 21552 36656 21560
tri 36656 21552 36664 21560 sw
rect 36532 21546 36664 21552
rect 36396 21544 36664 21546
tri 36664 21544 36672 21552 sw
rect 70802 21548 71000 21606
tri 36396 21536 36404 21544 ne
rect 36404 21536 36672 21544
tri 36672 21536 36680 21544 sw
tri 36404 21530 36410 21536 ne
rect 36410 21535 36680 21536
tri 36680 21535 36681 21536 sw
rect 36410 21530 36681 21535
tri 36410 21522 36418 21530 ne
rect 36418 21527 36681 21530
tri 36681 21527 36689 21535 sw
rect 36418 21522 36689 21527
tri 36418 21514 36426 21522 ne
rect 36426 21519 36689 21522
tri 36689 21519 36697 21527 sw
rect 36426 21514 36697 21519
tri 36426 21506 36434 21514 ne
rect 36434 21511 36697 21514
tri 36697 21511 36705 21519 sw
rect 36434 21506 36705 21511
tri 36434 21498 36442 21506 ne
rect 36442 21503 36705 21506
tri 36705 21503 36713 21511 sw
rect 36442 21498 36713 21503
tri 36442 21490 36450 21498 ne
rect 36450 21495 36713 21498
tri 36713 21495 36721 21503 sw
rect 70802 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
rect 36450 21490 36721 21495
tri 36450 21482 36458 21490 ne
rect 36458 21487 36721 21490
tri 36721 21487 36729 21495 sw
rect 36458 21482 36729 21487
tri 36458 21474 36466 21482 ne
rect 36466 21479 36729 21482
tri 36729 21479 36737 21487 sw
rect 36466 21474 36737 21479
tri 36466 21466 36474 21474 ne
rect 36474 21471 36737 21474
tri 36737 21471 36745 21479 sw
rect 36474 21466 36745 21471
tri 36474 21458 36482 21466 ne
rect 36482 21463 36745 21466
tri 36745 21463 36753 21471 sw
rect 36482 21460 36753 21463
rect 36482 21458 36618 21460
tri 36482 21450 36490 21458 ne
rect 36490 21450 36618 21458
tri 36490 21442 36498 21450 ne
rect 36498 21442 36618 21450
tri 36498 21434 36506 21442 ne
rect 36506 21434 36618 21442
tri 36506 21426 36514 21434 ne
rect 36514 21426 36618 21434
tri 36514 21418 36522 21426 ne
rect 36522 21418 36618 21426
tri 36522 21410 36530 21418 ne
rect 36530 21414 36618 21418
rect 36664 21455 36753 21460
tri 36753 21455 36761 21463 sw
rect 36664 21450 36761 21455
tri 36761 21450 36766 21455 sw
rect 36664 21442 36766 21450
tri 36766 21442 36774 21450 sw
rect 70802 21444 71000 21502
rect 36664 21434 36774 21442
tri 36774 21434 36782 21442 sw
rect 36664 21426 36782 21434
tri 36782 21426 36790 21434 sw
rect 36664 21418 36790 21426
tri 36790 21418 36798 21426 sw
rect 36664 21414 36798 21418
rect 36530 21410 36798 21414
tri 36798 21410 36806 21418 sw
tri 36530 21402 36538 21410 ne
rect 36538 21402 36806 21410
tri 36806 21402 36814 21410 sw
tri 36538 21394 36546 21402 ne
rect 36546 21394 36814 21402
tri 36814 21394 36822 21402 sw
rect 70802 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36546 21388 36552 21394 ne
rect 36552 21388 36822 21394
tri 36822 21388 36828 21394 sw
tri 36552 21380 36560 21388 ne
rect 36560 21380 36828 21388
tri 36828 21380 36836 21388 sw
tri 36560 21372 36568 21380 ne
rect 36568 21372 36836 21380
tri 36836 21372 36844 21380 sw
tri 36568 21364 36576 21372 ne
rect 36576 21364 36844 21372
tri 36844 21364 36852 21372 sw
tri 36576 21356 36584 21364 ne
rect 36584 21356 36852 21364
tri 36852 21356 36860 21364 sw
tri 36584 21348 36592 21356 ne
rect 36592 21348 36860 21356
tri 36860 21348 36868 21356 sw
tri 36592 21340 36600 21348 ne
rect 36600 21340 36868 21348
tri 36868 21340 36876 21348 sw
rect 70802 21340 71000 21398
tri 36600 21332 36608 21340 ne
rect 36608 21332 36876 21340
tri 36876 21332 36884 21340 sw
tri 36608 21324 36616 21332 ne
rect 36616 21328 36884 21332
rect 36616 21324 36750 21328
tri 36616 21316 36624 21324 ne
rect 36624 21316 36750 21324
tri 36624 21308 36632 21316 ne
rect 36632 21308 36750 21316
tri 36632 21300 36640 21308 ne
rect 36640 21300 36750 21308
tri 36640 21292 36648 21300 ne
rect 36648 21292 36750 21300
tri 36648 21284 36656 21292 ne
rect 36656 21284 36750 21292
tri 36656 21276 36664 21284 ne
rect 36664 21282 36750 21284
rect 36796 21324 36884 21328
tri 36884 21324 36892 21332 sw
rect 36796 21316 36892 21324
tri 36892 21316 36900 21324 sw
rect 36796 21308 36900 21316
tri 36900 21308 36908 21316 sw
rect 36796 21300 36908 21308
tri 36908 21300 36916 21308 sw
rect 36796 21292 36916 21300
tri 36916 21292 36924 21300 sw
rect 70802 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36796 21284 36924 21292
tri 36924 21284 36932 21292 sw
rect 36796 21282 36932 21284
rect 36664 21276 36932 21282
tri 36932 21276 36940 21284 sw
tri 36664 21268 36672 21276 ne
rect 36672 21271 36940 21276
tri 36940 21271 36945 21276 sw
rect 36672 21268 36945 21271
tri 36672 21260 36680 21268 ne
rect 36680 21263 36945 21268
tri 36945 21263 36953 21271 sw
rect 36680 21260 36953 21263
tri 36680 21252 36688 21260 ne
rect 36688 21255 36953 21260
tri 36953 21255 36961 21263 sw
rect 36688 21252 36961 21255
tri 36688 21251 36689 21252 ne
rect 36689 21251 36961 21252
tri 36689 21243 36697 21251 ne
rect 36697 21247 36961 21251
tri 36961 21247 36969 21255 sw
rect 36697 21243 36969 21247
tri 36697 21235 36705 21243 ne
rect 36705 21239 36969 21243
tri 36969 21239 36977 21247 sw
rect 36705 21235 36977 21239
tri 36705 21227 36713 21235 ne
rect 36713 21231 36977 21235
tri 36977 21231 36985 21239 sw
rect 70802 21236 71000 21294
rect 36713 21227 36985 21231
tri 36713 21219 36721 21227 ne
rect 36721 21223 36985 21227
tri 36985 21223 36993 21231 sw
rect 36721 21219 36993 21223
tri 36721 21211 36729 21219 ne
rect 36729 21215 36993 21219
tri 36993 21215 37001 21223 sw
rect 36729 21211 37001 21215
tri 36729 21203 36737 21211 ne
rect 36737 21207 37001 21211
tri 37001 21207 37009 21215 sw
rect 36737 21203 37009 21207
tri 36737 21195 36745 21203 ne
rect 36745 21199 37009 21203
tri 37009 21199 37017 21207 sw
rect 36745 21196 37017 21199
rect 36745 21195 36882 21196
tri 36745 21187 36753 21195 ne
rect 36753 21187 36882 21195
tri 36753 21179 36761 21187 ne
rect 36761 21179 36882 21187
tri 36761 21171 36769 21179 ne
rect 36769 21171 36882 21179
tri 36769 21163 36777 21171 ne
rect 36777 21163 36882 21171
tri 36777 21155 36785 21163 ne
rect 36785 21155 36882 21163
tri 36785 21147 36793 21155 ne
rect 36793 21150 36882 21155
rect 36928 21191 37017 21196
tri 37017 21191 37025 21199 sw
rect 36928 21187 37025 21191
tri 37025 21187 37029 21191 sw
rect 70802 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21179 37029 21187
tri 37029 21179 37037 21187 sw
rect 36928 21171 37037 21179
tri 37037 21171 37045 21179 sw
rect 36928 21163 37045 21171
tri 37045 21163 37053 21171 sw
rect 36928 21155 37053 21163
tri 37053 21155 37061 21163 sw
rect 36928 21150 37061 21155
rect 36793 21147 37061 21150
tri 37061 21147 37069 21155 sw
tri 36793 21139 36801 21147 ne
rect 36801 21139 37069 21147
tri 37069 21139 37077 21147 sw
tri 36801 21133 36807 21139 ne
rect 36807 21133 37077 21139
tri 36807 21125 36815 21133 ne
rect 36815 21131 37077 21133
tri 37077 21131 37085 21139 sw
rect 70802 21132 71000 21190
rect 36815 21125 37085 21131
tri 36815 21117 36823 21125 ne
rect 36823 21123 37085 21125
tri 37085 21123 37093 21131 sw
rect 36823 21117 37093 21123
tri 36823 21109 36831 21117 ne
rect 36831 21115 37093 21117
tri 37093 21115 37101 21123 sw
rect 36831 21109 37101 21115
tri 36831 21101 36839 21109 ne
rect 36839 21107 37101 21109
tri 37101 21107 37109 21115 sw
rect 36839 21101 37109 21107
tri 36839 21093 36847 21101 ne
rect 36847 21099 37109 21101
tri 37109 21099 37117 21107 sw
rect 36847 21093 37117 21099
tri 36847 21085 36855 21093 ne
rect 36855 21091 37117 21093
tri 37117 21091 37125 21099 sw
rect 36855 21085 37125 21091
tri 36855 21077 36863 21085 ne
rect 36863 21083 37125 21085
tri 37125 21083 37133 21091 sw
rect 70802 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 36863 21077 37133 21083
tri 36863 21069 36871 21077 ne
rect 36871 21075 37133 21077
tri 37133 21075 37141 21083 sw
rect 36871 21069 37141 21075
tri 36871 21061 36879 21069 ne
rect 36879 21067 37141 21069
tri 37141 21067 37149 21075 sw
rect 36879 21064 37149 21067
tri 37149 21064 37152 21067 sw
rect 36879 21061 37014 21064
tri 36879 21053 36887 21061 ne
rect 36887 21053 37014 21061
tri 36887 21045 36895 21053 ne
rect 36895 21045 37014 21053
tri 36895 21037 36903 21045 ne
rect 36903 21037 37014 21045
tri 36903 21029 36911 21037 ne
rect 36911 21029 37014 21037
tri 36911 21021 36919 21029 ne
rect 36919 21021 37014 21029
tri 36919 21015 36925 21021 ne
rect 36925 21018 37014 21021
rect 37060 21056 37152 21064
tri 37152 21056 37160 21064 sw
rect 37060 21048 37160 21056
tri 37160 21048 37168 21056 sw
rect 37060 21040 37168 21048
tri 37168 21040 37176 21048 sw
rect 37060 21032 37176 21040
tri 37176 21032 37184 21040 sw
rect 37060 21024 37184 21032
tri 37184 21024 37192 21032 sw
rect 70802 21028 71000 21086
rect 37060 21018 37192 21024
rect 36925 21016 37192 21018
tri 37192 21016 37200 21024 sw
rect 36925 21015 37200 21016
tri 36925 21007 36933 21015 ne
rect 36933 21008 37200 21015
tri 37200 21008 37208 21016 sw
rect 36933 21007 37208 21008
tri 36933 20999 36941 21007 ne
rect 36941 21000 37208 21007
tri 37208 21000 37216 21008 sw
rect 36941 20999 37216 21000
tri 36941 20991 36949 20999 ne
rect 36949 20992 37216 20999
tri 37216 20992 37224 21000 sw
rect 36949 20991 37224 20992
tri 36949 20983 36957 20991 ne
rect 36957 20984 37224 20991
tri 37224 20984 37232 20992 sw
rect 36957 20983 37232 20984
tri 36957 20975 36965 20983 ne
rect 36965 20976 37232 20983
tri 37232 20976 37240 20984 sw
rect 70802 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
rect 36965 20975 37240 20976
tri 36965 20967 36973 20975 ne
rect 36973 20968 37240 20975
tri 37240 20968 37248 20976 sw
rect 36973 20967 37248 20968
tri 36973 20959 36981 20967 ne
rect 36981 20960 37248 20967
tri 37248 20960 37256 20968 sw
rect 36981 20959 37256 20960
tri 36981 20951 36989 20959 ne
rect 36989 20952 37256 20959
tri 37256 20952 37264 20960 sw
rect 36989 20951 37264 20952
tri 37264 20951 37265 20952 sw
tri 36989 20943 36997 20951 ne
rect 36997 20943 37265 20951
tri 37265 20943 37273 20951 sw
tri 36997 20935 37005 20943 ne
rect 37005 20935 37273 20943
tri 37273 20935 37281 20943 sw
tri 37005 20931 37009 20935 ne
rect 37009 20932 37281 20935
rect 37009 20931 37146 20932
tri 37009 20927 37013 20931 ne
rect 37013 20927 37146 20931
tri 37013 20919 37021 20927 ne
rect 37021 20919 37146 20927
tri 37021 20911 37029 20919 ne
rect 37029 20911 37146 20919
tri 37029 20903 37037 20911 ne
rect 37037 20903 37146 20911
tri 37037 20895 37045 20903 ne
rect 37045 20895 37146 20903
tri 37045 20887 37053 20895 ne
rect 37053 20887 37146 20895
tri 37053 20879 37061 20887 ne
rect 37061 20886 37146 20887
rect 37192 20927 37281 20932
tri 37281 20927 37289 20935 sw
rect 37192 20919 37289 20927
tri 37289 20919 37297 20927 sw
rect 70802 20924 71000 20982
rect 37192 20911 37297 20919
tri 37297 20911 37305 20919 sw
rect 37192 20903 37305 20911
tri 37305 20903 37313 20911 sw
rect 37192 20895 37313 20903
tri 37313 20895 37321 20903 sw
rect 37192 20887 37321 20895
tri 37321 20887 37329 20895 sw
rect 37192 20886 37329 20887
rect 37061 20879 37329 20886
tri 37329 20879 37337 20887 sw
tri 37061 20871 37069 20879 ne
rect 37069 20873 37337 20879
tri 37337 20873 37343 20879 sw
rect 70802 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 37069 20871 37343 20873
tri 37069 20863 37077 20871 ne
rect 37077 20865 37343 20871
tri 37343 20865 37351 20873 sw
rect 37077 20863 37351 20865
tri 37077 20860 37080 20863 ne
rect 37080 20860 37351 20863
tri 37080 20852 37088 20860 ne
rect 37088 20857 37351 20860
tri 37351 20857 37359 20865 sw
rect 37088 20852 37359 20857
tri 37088 20844 37096 20852 ne
rect 37096 20849 37359 20852
tri 37359 20849 37367 20857 sw
rect 37096 20844 37367 20849
tri 37096 20836 37104 20844 ne
rect 37104 20841 37367 20844
tri 37367 20841 37375 20849 sw
rect 37104 20836 37375 20841
tri 37104 20828 37112 20836 ne
rect 37112 20833 37375 20836
tri 37375 20833 37383 20841 sw
rect 37112 20828 37383 20833
tri 37112 20820 37120 20828 ne
rect 37120 20825 37383 20828
tri 37383 20825 37391 20833 sw
rect 37120 20820 37391 20825
tri 37120 20812 37128 20820 ne
rect 37128 20817 37391 20820
tri 37391 20817 37399 20825 sw
rect 70802 20820 71000 20878
rect 37128 20812 37399 20817
tri 37128 20804 37136 20812 ne
rect 37136 20809 37399 20812
tri 37399 20809 37407 20817 sw
rect 37136 20804 37407 20809
tri 37136 20796 37144 20804 ne
rect 37144 20801 37407 20804
tri 37407 20801 37415 20809 sw
rect 37144 20800 37415 20801
rect 37144 20796 37278 20800
tri 37144 20788 37152 20796 ne
rect 37152 20788 37278 20796
tri 37152 20780 37160 20788 ne
rect 37160 20780 37278 20788
tri 37160 20772 37168 20780 ne
rect 37168 20772 37278 20780
tri 37168 20764 37176 20772 ne
rect 37176 20764 37278 20772
tri 37176 20756 37184 20764 ne
rect 37184 20756 37278 20764
tri 37184 20748 37192 20756 ne
rect 37192 20754 37278 20756
rect 37324 20793 37415 20800
tri 37415 20793 37423 20801 sw
rect 37324 20785 37423 20793
tri 37423 20785 37431 20793 sw
rect 37324 20777 37431 20785
tri 37431 20777 37439 20785 sw
rect 37324 20769 37439 20777
tri 37439 20769 37447 20777 sw
rect 70802 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 37324 20761 37447 20769
tri 37447 20761 37455 20769 sw
rect 37324 20754 37455 20761
rect 37192 20753 37455 20754
tri 37455 20753 37463 20761 sw
rect 37192 20748 37463 20753
tri 37192 20740 37200 20748 ne
rect 37200 20745 37463 20748
tri 37463 20745 37471 20753 sw
rect 37200 20740 37471 20745
tri 37200 20732 37208 20740 ne
rect 37208 20739 37471 20740
tri 37471 20739 37477 20745 sw
rect 37208 20732 37477 20739
tri 37208 20724 37216 20732 ne
rect 37216 20731 37477 20732
tri 37477 20731 37485 20739 sw
rect 37216 20724 37485 20731
tri 37216 20723 37217 20724 ne
rect 37217 20723 37485 20724
tri 37485 20723 37493 20731 sw
tri 37217 20715 37225 20723 ne
rect 37225 20715 37493 20723
tri 37493 20715 37501 20723 sw
rect 70802 20716 71000 20774
tri 37225 20707 37233 20715 ne
rect 37233 20707 37501 20715
tri 37501 20707 37509 20715 sw
tri 37233 20699 37241 20707 ne
rect 37241 20699 37509 20707
tri 37509 20699 37517 20707 sw
tri 37241 20691 37249 20699 ne
rect 37249 20691 37517 20699
tri 37517 20691 37525 20699 sw
tri 37249 20683 37257 20691 ne
rect 37257 20683 37525 20691
tri 37525 20683 37533 20691 sw
tri 37257 20675 37265 20683 ne
rect 37265 20675 37533 20683
tri 37533 20675 37541 20683 sw
tri 37265 20667 37273 20675 ne
rect 37273 20668 37541 20675
rect 37273 20667 37410 20668
tri 37273 20659 37281 20667 ne
rect 37281 20659 37410 20667
tri 37281 20651 37289 20659 ne
rect 37289 20651 37410 20659
tri 37289 20643 37297 20651 ne
rect 37297 20643 37410 20651
tri 37297 20635 37305 20643 ne
rect 37305 20635 37410 20643
tri 37305 20627 37313 20635 ne
rect 37313 20627 37410 20635
tri 37313 20619 37321 20627 ne
rect 37321 20622 37410 20627
rect 37456 20667 37541 20668
tri 37541 20667 37549 20675 sw
rect 70802 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 37456 20659 37549 20667
tri 37549 20659 37557 20667 sw
rect 37456 20651 37557 20659
tri 37557 20651 37565 20659 sw
rect 37456 20643 37565 20651
tri 37565 20643 37573 20651 sw
rect 37456 20635 37573 20643
tri 37573 20635 37581 20643 sw
rect 37456 20627 37581 20635
tri 37581 20627 37589 20635 sw
rect 37456 20622 37589 20627
rect 37321 20619 37589 20622
tri 37589 20619 37597 20627 sw
tri 37321 20611 37329 20619 ne
rect 37329 20611 37597 20619
tri 37597 20611 37605 20619 sw
rect 70802 20612 71000 20670
tri 37329 20603 37337 20611 ne
rect 37337 20603 37605 20611
tri 37605 20603 37613 20611 sw
tri 37337 20597 37343 20603 ne
rect 37343 20597 37613 20603
tri 37613 20597 37619 20603 sw
tri 37343 20589 37351 20597 ne
rect 37351 20589 37619 20597
tri 37619 20589 37627 20597 sw
tri 37351 20581 37359 20589 ne
rect 37359 20581 37627 20589
tri 37627 20581 37635 20589 sw
tri 37359 20573 37367 20581 ne
rect 37367 20573 37635 20581
tri 37635 20573 37643 20581 sw
tri 37367 20565 37375 20573 ne
rect 37375 20565 37643 20573
tri 37643 20565 37651 20573 sw
rect 70802 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
tri 37375 20557 37383 20565 ne
rect 37383 20557 37651 20565
tri 37651 20557 37659 20565 sw
tri 37383 20549 37391 20557 ne
rect 37391 20549 37659 20557
tri 37659 20549 37667 20557 sw
tri 37391 20541 37399 20549 ne
rect 37399 20541 37667 20549
tri 37667 20541 37675 20549 sw
tri 37399 20533 37407 20541 ne
rect 37407 20536 37675 20541
rect 37407 20533 37542 20536
tri 37407 20525 37415 20533 ne
rect 37415 20525 37542 20533
tri 37415 20517 37423 20525 ne
rect 37423 20517 37542 20525
tri 37423 20509 37431 20517 ne
rect 37431 20509 37542 20517
tri 37431 20501 37439 20509 ne
rect 37439 20501 37542 20509
tri 37439 20493 37447 20501 ne
rect 37447 20493 37542 20501
tri 37447 20485 37455 20493 ne
rect 37455 20490 37542 20493
rect 37588 20533 37675 20536
tri 37675 20533 37683 20541 sw
rect 37588 20525 37683 20533
tri 37683 20525 37691 20533 sw
rect 37588 20517 37691 20525
tri 37691 20517 37699 20525 sw
rect 37588 20509 37699 20517
tri 37699 20509 37707 20517 sw
rect 37588 20501 37707 20509
tri 37707 20501 37715 20509 sw
rect 70802 20508 71000 20566
rect 37588 20493 37715 20501
tri 37715 20493 37723 20501 sw
rect 37588 20490 37723 20493
rect 37455 20487 37723 20490
tri 37723 20487 37729 20493 sw
rect 37455 20485 37729 20487
tri 37455 20477 37463 20485 ne
rect 37463 20479 37729 20485
tri 37729 20479 37737 20487 sw
rect 37463 20477 37737 20479
tri 37463 20474 37466 20477 ne
rect 37466 20474 37737 20477
tri 37466 20466 37474 20474 ne
rect 37474 20471 37737 20474
tri 37737 20471 37745 20479 sw
rect 37474 20466 37745 20471
tri 37474 20458 37482 20466 ne
rect 37482 20463 37745 20466
tri 37745 20463 37753 20471 sw
rect 37482 20458 37753 20463
tri 37482 20450 37490 20458 ne
rect 37490 20455 37753 20458
tri 37753 20455 37761 20463 sw
rect 70802 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
rect 37490 20450 37761 20455
tri 37490 20442 37498 20450 ne
rect 37498 20447 37761 20450
tri 37761 20447 37769 20455 sw
rect 37498 20442 37769 20447
tri 37498 20434 37506 20442 ne
rect 37506 20439 37769 20442
tri 37769 20439 37777 20447 sw
rect 37506 20434 37777 20439
tri 37506 20426 37514 20434 ne
rect 37514 20431 37777 20434
tri 37777 20431 37785 20439 sw
rect 37514 20426 37785 20431
tri 37514 20418 37522 20426 ne
rect 37522 20423 37785 20426
tri 37785 20423 37793 20431 sw
rect 37522 20418 37793 20423
tri 37522 20410 37530 20418 ne
rect 37530 20415 37793 20418
tri 37793 20415 37801 20423 sw
rect 37530 20410 37801 20415
tri 37530 20402 37538 20410 ne
rect 37538 20407 37801 20410
tri 37801 20407 37809 20415 sw
rect 37538 20404 37809 20407
rect 37538 20402 37674 20404
tri 37538 20394 37546 20402 ne
rect 37546 20394 37674 20402
tri 37546 20386 37554 20394 ne
rect 37554 20386 37674 20394
tri 37554 20378 37562 20386 ne
rect 37562 20378 37674 20386
tri 37562 20370 37570 20378 ne
rect 37570 20370 37674 20378
tri 37570 20362 37578 20370 ne
rect 37578 20362 37674 20370
tri 37578 20354 37586 20362 ne
rect 37586 20358 37674 20362
rect 37720 20402 37809 20404
tri 37809 20402 37814 20407 sw
rect 70802 20404 71000 20462
rect 37720 20394 37814 20402
tri 37814 20394 37822 20402 sw
rect 37720 20386 37822 20394
tri 37822 20386 37830 20394 sw
rect 37720 20378 37830 20386
tri 37830 20378 37838 20386 sw
rect 37720 20370 37838 20378
tri 37838 20370 37846 20378 sw
rect 37720 20362 37846 20370
tri 37846 20362 37854 20370 sw
rect 37720 20358 37854 20362
rect 37586 20354 37854 20358
tri 37854 20354 37862 20362 sw
rect 70802 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37586 20346 37594 20354 ne
rect 37594 20346 37862 20354
tri 37862 20346 37870 20354 sw
tri 37594 20338 37602 20346 ne
rect 37602 20338 37870 20346
tri 37870 20338 37878 20346 sw
tri 37602 20330 37610 20338 ne
rect 37610 20337 37878 20338
tri 37878 20337 37879 20338 sw
rect 37610 20330 37879 20337
tri 37610 20329 37611 20330 ne
rect 37611 20329 37879 20330
tri 37879 20329 37887 20337 sw
tri 37611 20321 37619 20329 ne
rect 37619 20321 37887 20329
tri 37887 20321 37895 20329 sw
tri 37619 20313 37627 20321 ne
rect 37627 20313 37895 20321
tri 37895 20313 37903 20321 sw
tri 37627 20305 37635 20313 ne
rect 37635 20305 37903 20313
tri 37903 20305 37911 20313 sw
tri 37635 20297 37643 20305 ne
rect 37643 20297 37911 20305
tri 37911 20297 37919 20305 sw
rect 70802 20300 71000 20358
tri 37643 20289 37651 20297 ne
rect 37651 20289 37919 20297
tri 37919 20289 37927 20297 sw
tri 37651 20281 37659 20289 ne
rect 37659 20281 37927 20289
tri 37927 20281 37935 20289 sw
tri 37659 20273 37667 20281 ne
rect 37667 20273 37935 20281
tri 37935 20273 37943 20281 sw
tri 37667 20265 37675 20273 ne
rect 37675 20272 37943 20273
rect 37675 20265 37806 20272
tri 37675 20257 37683 20265 ne
rect 37683 20257 37806 20265
tri 37683 20249 37691 20257 ne
rect 37691 20249 37806 20257
tri 37691 20241 37699 20249 ne
rect 37699 20241 37806 20249
tri 37699 20233 37707 20241 ne
rect 37707 20233 37806 20241
tri 37707 20225 37715 20233 ne
rect 37715 20226 37806 20233
rect 37852 20265 37943 20272
tri 37943 20265 37951 20273 sw
rect 37852 20257 37951 20265
tri 37951 20257 37959 20265 sw
rect 37852 20249 37959 20257
tri 37959 20249 37967 20257 sw
rect 70802 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20241 37967 20249
tri 37967 20241 37975 20249 sw
rect 37852 20233 37975 20241
tri 37975 20233 37983 20241 sw
rect 37852 20226 37983 20233
rect 37715 20225 37983 20226
tri 37983 20225 37991 20233 sw
tri 37715 20217 37723 20225 ne
rect 37723 20217 37991 20225
tri 37991 20217 37999 20225 sw
tri 37723 20209 37731 20217 ne
rect 37731 20209 37999 20217
tri 37999 20209 38007 20217 sw
tri 37731 20203 37737 20209 ne
rect 37737 20203 38007 20209
tri 38007 20203 38013 20209 sw
tri 37737 20195 37745 20203 ne
rect 37745 20195 38013 20203
tri 38013 20195 38021 20203 sw
rect 70802 20196 71000 20254
tri 37745 20187 37753 20195 ne
rect 37753 20187 38021 20195
tri 38021 20187 38029 20195 sw
tri 37753 20179 37761 20187 ne
rect 37761 20179 38029 20187
tri 38029 20179 38037 20187 sw
tri 37761 20171 37769 20179 ne
rect 37769 20171 38037 20179
tri 38037 20171 38045 20179 sw
tri 37769 20163 37777 20171 ne
rect 37777 20163 38045 20171
tri 38045 20163 38053 20171 sw
tri 37777 20155 37785 20163 ne
rect 37785 20155 38053 20163
tri 38053 20155 38061 20163 sw
tri 37785 20147 37793 20155 ne
rect 37793 20147 38061 20155
tri 38061 20147 38069 20155 sw
rect 70802 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
tri 37793 20139 37801 20147 ne
rect 37801 20140 38069 20147
rect 37801 20139 37938 20140
tri 37801 20131 37809 20139 ne
rect 37809 20131 37938 20139
tri 37809 20123 37817 20131 ne
rect 37817 20123 37938 20131
tri 37817 20115 37825 20123 ne
rect 37825 20115 37938 20123
tri 37825 20107 37833 20115 ne
rect 37833 20107 37938 20115
tri 37833 20099 37841 20107 ne
rect 37841 20099 37938 20107
tri 37841 20091 37849 20099 ne
rect 37849 20094 37938 20099
rect 37984 20139 38069 20140
tri 38069 20139 38077 20147 sw
rect 37984 20131 38077 20139
tri 38077 20131 38085 20139 sw
rect 37984 20123 38085 20131
tri 38085 20123 38093 20131 sw
rect 37984 20115 38093 20123
tri 38093 20115 38101 20123 sw
rect 37984 20107 38101 20115
tri 38101 20107 38109 20115 sw
rect 37984 20099 38109 20107
tri 38109 20099 38117 20107 sw
rect 37984 20094 38117 20099
rect 37849 20091 38117 20094
tri 38117 20091 38125 20099 sw
rect 70802 20092 71000 20150
tri 37849 20083 37857 20091 ne
rect 37857 20083 38125 20091
tri 38125 20083 38133 20091 sw
tri 37857 20075 37865 20083 ne
rect 37865 20075 38133 20083
tri 38133 20075 38141 20083 sw
tri 37865 20067 37873 20075 ne
rect 37873 20067 38141 20075
tri 38141 20067 38149 20075 sw
tri 37873 20066 37874 20067 ne
rect 37874 20066 38149 20067
tri 37874 20058 37882 20066 ne
rect 37882 20059 38149 20066
tri 38149 20059 38157 20067 sw
rect 37882 20058 38157 20059
tri 37882 20050 37890 20058 ne
rect 37890 20051 38157 20058
tri 38157 20051 38165 20059 sw
rect 37890 20050 38165 20051
tri 37890 20042 37898 20050 ne
rect 37898 20043 38165 20050
tri 38165 20043 38173 20051 sw
rect 70802 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
rect 37898 20042 38173 20043
tri 37898 20034 37906 20042 ne
rect 37906 20035 38173 20042
tri 38173 20035 38181 20043 sw
rect 37906 20034 38181 20035
tri 37906 20026 37914 20034 ne
rect 37914 20027 38181 20034
tri 38181 20027 38189 20035 sw
rect 37914 20026 38189 20027
tri 37914 20018 37922 20026 ne
rect 37922 20019 38189 20026
tri 38189 20019 38197 20027 sw
rect 37922 20018 38197 20019
tri 37922 20010 37930 20018 ne
rect 37930 20011 38197 20018
tri 38197 20011 38205 20019 sw
rect 37930 20010 38205 20011
tri 37930 20002 37938 20010 ne
rect 37938 20008 38205 20010
rect 37938 20002 38070 20008
tri 37938 19994 37946 20002 ne
rect 37946 19994 38070 20002
tri 37946 19986 37954 19994 ne
rect 37954 19986 38070 19994
tri 37954 19978 37962 19986 ne
rect 37962 19978 38070 19986
tri 37962 19970 37970 19978 ne
rect 37970 19970 38070 19978
tri 37970 19962 37978 19970 ne
rect 37978 19962 38070 19970
rect 38116 20003 38205 20008
tri 38205 20003 38213 20011 sw
rect 38116 19995 38213 20003
tri 38213 19995 38221 20003 sw
rect 38116 19987 38221 19995
tri 38221 19987 38229 19995 sw
rect 70802 19988 71000 20046
rect 38116 19979 38229 19987
tri 38229 19979 38237 19987 sw
rect 38116 19971 38237 19979
tri 38237 19971 38245 19979 sw
rect 38116 19963 38245 19971
tri 38245 19963 38253 19971 sw
rect 38116 19962 38253 19963
tri 37978 19954 37986 19962 ne
rect 37986 19955 38253 19962
tri 38253 19955 38261 19963 sw
rect 37986 19954 38261 19955
tri 37986 19946 37994 19954 ne
rect 37994 19948 38261 19954
tri 38261 19948 38268 19955 sw
rect 37994 19946 38268 19948
tri 37994 19938 38002 19946 ne
rect 38002 19940 38268 19946
tri 38268 19940 38276 19948 sw
rect 70802 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 38002 19938 38276 19940
tri 38002 19930 38010 19938 ne
rect 38010 19932 38276 19938
tri 38276 19932 38284 19940 sw
rect 38010 19930 38284 19932
tri 38010 19922 38018 19930 ne
rect 38018 19924 38284 19930
tri 38284 19924 38292 19932 sw
rect 38018 19922 38292 19924
tri 38018 19914 38026 19922 ne
rect 38026 19916 38292 19922
tri 38292 19916 38300 19924 sw
rect 38026 19914 38300 19916
tri 38026 19906 38034 19914 ne
rect 38034 19908 38300 19914
tri 38300 19908 38308 19916 sw
rect 38034 19906 38308 19908
tri 38034 19898 38042 19906 ne
rect 38042 19900 38308 19906
tri 38308 19900 38316 19908 sw
rect 38042 19898 38316 19900
tri 38042 19890 38050 19898 ne
rect 38050 19892 38316 19898
tri 38316 19892 38324 19900 sw
rect 38050 19890 38324 19892
tri 38050 19882 38058 19890 ne
rect 38058 19884 38324 19890
tri 38324 19884 38332 19892 sw
rect 70802 19884 71000 19942
rect 38058 19882 38332 19884
tri 38058 19874 38066 19882 ne
rect 38066 19876 38332 19882
tri 38332 19876 38340 19884 sw
rect 38066 19874 38202 19876
tri 38066 19870 38070 19874 ne
rect 38070 19870 38202 19874
tri 38070 19866 38074 19870 ne
rect 38074 19866 38202 19870
tri 38074 19858 38082 19866 ne
rect 38082 19858 38202 19866
tri 38082 19850 38090 19858 ne
rect 38090 19850 38202 19858
tri 38090 19842 38098 19850 ne
rect 38098 19842 38202 19850
tri 38098 19834 38106 19842 ne
rect 38106 19834 38202 19842
tri 38106 19826 38114 19834 ne
rect 38114 19830 38202 19834
rect 38248 19868 38340 19876
tri 38340 19868 38348 19876 sw
rect 38248 19860 38348 19868
tri 38348 19860 38356 19868 sw
rect 38248 19852 38356 19860
tri 38356 19852 38364 19860 sw
rect 38248 19844 38364 19852
tri 38364 19844 38372 19852 sw
rect 38248 19836 38372 19844
tri 38372 19836 38380 19844 sw
rect 70802 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 38248 19830 38380 19836
rect 38114 19828 38380 19830
tri 38380 19828 38388 19836 sw
rect 38114 19826 38388 19828
tri 38114 19818 38122 19826 ne
rect 38122 19820 38388 19826
tri 38388 19820 38396 19828 sw
rect 38122 19818 38396 19820
tri 38122 19810 38130 19818 ne
rect 38130 19812 38396 19818
tri 38396 19812 38404 19820 sw
rect 38130 19810 38404 19812
tri 38130 19802 38138 19810 ne
rect 38138 19804 38404 19810
tri 38404 19804 38412 19812 sw
rect 38138 19802 38412 19804
tri 38138 19794 38146 19802 ne
rect 38146 19796 38412 19802
tri 38412 19796 38420 19804 sw
rect 38146 19794 38420 19796
tri 38146 19786 38154 19794 ne
rect 38154 19788 38420 19794
tri 38420 19788 38428 19796 sw
rect 38154 19786 38428 19788
tri 38154 19778 38162 19786 ne
rect 38162 19780 38428 19786
tri 38428 19780 38436 19788 sw
rect 70802 19780 71000 19838
rect 38162 19778 38436 19780
tri 38162 19770 38170 19778 ne
rect 38170 19772 38436 19778
tri 38436 19772 38444 19780 sw
rect 38170 19770 38444 19772
tri 38170 19762 38178 19770 ne
rect 38178 19765 38444 19770
tri 38444 19765 38451 19772 sw
rect 38178 19762 38451 19765
tri 38178 19754 38186 19762 ne
rect 38186 19757 38451 19762
tri 38451 19757 38459 19765 sw
rect 38186 19754 38459 19757
tri 38186 19746 38194 19754 ne
rect 38194 19749 38459 19754
tri 38459 19749 38467 19757 sw
rect 38194 19746 38467 19749
tri 38194 19738 38202 19746 ne
rect 38202 19744 38467 19746
rect 38202 19738 38334 19744
tri 38202 19732 38208 19738 ne
rect 38208 19732 38334 19738
tri 38208 19724 38216 19732 ne
rect 38216 19724 38334 19732
tri 38216 19716 38224 19724 ne
rect 38224 19716 38334 19724
tri 38224 19708 38232 19716 ne
rect 38232 19708 38334 19716
tri 38232 19700 38240 19708 ne
rect 38240 19700 38334 19708
tri 38240 19692 38248 19700 ne
rect 38248 19698 38334 19700
rect 38380 19741 38467 19744
tri 38467 19741 38475 19749 sw
rect 38380 19733 38475 19741
tri 38475 19733 38483 19741 sw
rect 70802 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 38380 19725 38483 19733
tri 38483 19725 38491 19733 sw
rect 38380 19717 38491 19725
tri 38491 19717 38499 19725 sw
rect 38380 19709 38499 19717
tri 38499 19709 38507 19717 sw
rect 38380 19701 38507 19709
tri 38507 19701 38515 19709 sw
rect 38380 19698 38515 19701
rect 38248 19693 38515 19698
tri 38515 19693 38523 19701 sw
rect 38248 19692 38523 19693
tri 38248 19684 38256 19692 ne
rect 38256 19685 38523 19692
tri 38523 19685 38531 19693 sw
rect 38256 19684 38531 19685
tri 38256 19676 38264 19684 ne
rect 38264 19677 38531 19684
tri 38531 19677 38539 19685 sw
rect 38264 19676 38539 19677
tri 38264 19668 38272 19676 ne
rect 38272 19669 38539 19676
tri 38539 19669 38547 19677 sw
rect 70802 19676 71000 19734
rect 38272 19668 38547 19669
tri 38272 19660 38280 19668 ne
rect 38280 19661 38547 19668
tri 38547 19661 38555 19669 sw
rect 38280 19660 38555 19661
tri 38280 19652 38288 19660 ne
rect 38288 19653 38555 19660
tri 38555 19653 38563 19661 sw
rect 38288 19652 38563 19653
tri 38288 19644 38296 19652 ne
rect 38296 19645 38563 19652
tri 38563 19645 38571 19653 sw
rect 38296 19644 38571 19645
tri 38296 19636 38304 19644 ne
rect 38304 19637 38571 19644
tri 38571 19637 38579 19645 sw
rect 38304 19636 38579 19637
tri 38304 19628 38312 19636 ne
rect 38312 19635 38579 19636
tri 38579 19635 38581 19637 sw
rect 38312 19628 38581 19635
tri 38312 19620 38320 19628 ne
rect 38320 19627 38581 19628
tri 38581 19627 38589 19635 sw
rect 70802 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38320 19620 38589 19627
tri 38320 19612 38328 19620 ne
rect 38328 19619 38589 19620
tri 38589 19619 38597 19627 sw
rect 38328 19612 38597 19619
tri 38328 19608 38332 19612 ne
rect 38332 19608 38466 19612
tri 38332 19604 38336 19608 ne
rect 38336 19604 38466 19608
tri 38336 19596 38344 19604 ne
rect 38344 19596 38466 19604
tri 38344 19588 38352 19596 ne
rect 38352 19588 38466 19596
tri 38352 19580 38360 19588 ne
rect 38360 19580 38466 19588
tri 38360 19572 38368 19580 ne
rect 38368 19572 38466 19580
tri 38368 19564 38376 19572 ne
rect 38376 19566 38466 19572
rect 38512 19611 38597 19612
tri 38597 19611 38605 19619 sw
rect 38512 19603 38605 19611
tri 38605 19603 38613 19611 sw
rect 38512 19595 38613 19603
tri 38613 19595 38621 19603 sw
rect 38512 19587 38621 19595
tri 38621 19587 38629 19595 sw
rect 38512 19579 38629 19587
tri 38629 19579 38637 19587 sw
rect 38512 19571 38637 19579
tri 38637 19571 38645 19579 sw
rect 70802 19572 71000 19630
rect 38512 19566 38645 19571
rect 38376 19564 38645 19566
tri 38376 19556 38384 19564 ne
rect 38384 19563 38645 19564
tri 38645 19563 38653 19571 sw
rect 38384 19556 38653 19563
tri 38384 19548 38392 19556 ne
rect 38392 19555 38653 19556
tri 38653 19555 38661 19563 sw
rect 38392 19548 38661 19555
tri 38392 19540 38400 19548 ne
rect 38400 19547 38661 19548
tri 38661 19547 38669 19555 sw
rect 38400 19546 38669 19547
tri 38669 19546 38670 19547 sw
rect 38400 19540 38670 19546
tri 38400 19538 38402 19540 ne
rect 38402 19538 38670 19540
tri 38670 19538 38678 19546 sw
tri 38402 19530 38410 19538 ne
rect 38410 19530 38678 19538
tri 38678 19530 38686 19538 sw
tri 38410 19522 38418 19530 ne
rect 38418 19522 38686 19530
tri 38686 19522 38694 19530 sw
rect 70802 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38418 19514 38426 19522 ne
rect 38426 19514 38694 19522
tri 38694 19514 38702 19522 sw
tri 38426 19506 38434 19514 ne
rect 38434 19506 38702 19514
tri 38702 19506 38710 19514 sw
tri 38434 19498 38442 19506 ne
rect 38442 19498 38710 19506
tri 38710 19498 38718 19506 sw
tri 38442 19490 38450 19498 ne
rect 38450 19490 38718 19498
tri 38718 19490 38726 19498 sw
tri 38450 19482 38458 19490 ne
rect 38458 19482 38726 19490
tri 38726 19482 38734 19490 sw
tri 38458 19474 38466 19482 ne
rect 38466 19480 38734 19482
rect 38466 19474 38598 19480
tri 38466 19466 38474 19474 ne
rect 38474 19466 38598 19474
tri 38474 19458 38482 19466 ne
rect 38482 19458 38598 19466
tri 38482 19450 38490 19458 ne
rect 38490 19450 38598 19458
tri 38490 19442 38498 19450 ne
rect 38498 19442 38598 19450
tri 38498 19434 38506 19442 ne
rect 38506 19434 38598 19442
rect 38644 19474 38734 19480
tri 38734 19474 38742 19482 sw
rect 38644 19466 38742 19474
tri 38742 19466 38750 19474 sw
rect 70802 19468 71000 19526
rect 38644 19458 38750 19466
tri 38750 19458 38758 19466 sw
rect 38644 19450 38758 19458
tri 38758 19450 38766 19458 sw
rect 38644 19442 38766 19450
tri 38766 19442 38774 19450 sw
rect 38644 19437 38774 19442
tri 38774 19437 38779 19442 sw
rect 38644 19434 38779 19437
tri 38506 19426 38514 19434 ne
rect 38514 19429 38779 19434
tri 38779 19429 38787 19437 sw
rect 38514 19426 38787 19429
tri 38514 19418 38522 19426 ne
rect 38522 19421 38787 19426
tri 38787 19421 38795 19429 sw
rect 70802 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
rect 38522 19418 38795 19421
tri 38522 19415 38525 19418 ne
rect 38525 19415 38795 19418
tri 38525 19407 38533 19415 ne
rect 38533 19413 38795 19415
tri 38795 19413 38803 19421 sw
rect 38533 19407 38803 19413
tri 38533 19399 38541 19407 ne
rect 38541 19405 38803 19407
tri 38803 19405 38811 19413 sw
rect 38541 19399 38811 19405
tri 38541 19391 38549 19399 ne
rect 38549 19397 38811 19399
tri 38811 19397 38819 19405 sw
rect 38549 19391 38819 19397
tri 38549 19383 38557 19391 ne
rect 38557 19389 38819 19391
tri 38819 19389 38827 19397 sw
rect 38557 19383 38827 19389
tri 38557 19375 38565 19383 ne
rect 38565 19381 38827 19383
tri 38827 19381 38835 19389 sw
rect 38565 19377 38835 19381
tri 38835 19377 38839 19381 sw
rect 38565 19375 38839 19377
tri 38565 19367 38573 19375 ne
rect 38573 19373 38839 19375
tri 38839 19373 38843 19377 sw
rect 38573 19367 38843 19373
tri 38573 19359 38581 19367 ne
rect 38581 19365 38843 19367
tri 38843 19365 38851 19373 sw
rect 38581 19359 38851 19365
tri 38851 19359 38857 19365 sw
rect 70802 19364 71000 19422
tri 38581 19355 38585 19359 ne
rect 38585 19355 38857 19359
tri 38585 19351 38589 19355 ne
rect 38589 19351 38857 19355
tri 38857 19351 38865 19359 sw
tri 38589 19343 38597 19351 ne
rect 38597 19348 38865 19351
rect 38597 19343 38730 19348
tri 38597 19335 38605 19343 ne
rect 38605 19335 38730 19343
tri 38605 19327 38613 19335 ne
rect 38613 19327 38730 19335
tri 38613 19319 38621 19327 ne
rect 38621 19319 38730 19327
tri 38621 19311 38629 19319 ne
rect 38629 19311 38730 19319
tri 38629 19303 38637 19311 ne
rect 38637 19303 38730 19311
tri 38637 19295 38645 19303 ne
rect 38645 19302 38730 19303
rect 38776 19343 38865 19348
tri 38865 19343 38873 19351 sw
rect 38776 19335 38873 19343
tri 38873 19335 38881 19343 sw
rect 38776 19327 38881 19335
tri 38881 19327 38889 19335 sw
rect 38776 19319 38889 19327
tri 38889 19319 38897 19327 sw
rect 38776 19311 38897 19319
tri 38897 19311 38905 19319 sw
rect 70802 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 38776 19303 38905 19311
tri 38905 19303 38913 19311 sw
rect 38776 19302 38913 19303
rect 38645 19298 38913 19302
tri 38913 19298 38918 19303 sw
rect 38645 19295 38918 19298
tri 38645 19287 38653 19295 ne
rect 38653 19290 38918 19295
tri 38918 19290 38926 19298 sw
rect 38653 19287 38926 19290
tri 38653 19279 38661 19287 ne
rect 38661 19282 38926 19287
tri 38926 19282 38934 19290 sw
rect 38661 19279 38934 19282
tri 38661 19274 38666 19279 ne
rect 38666 19274 38934 19279
tri 38934 19274 38942 19282 sw
tri 38666 19266 38674 19274 ne
rect 38674 19266 38942 19274
tri 38942 19266 38950 19274 sw
tri 38674 19258 38682 19266 ne
rect 38682 19258 38950 19266
tri 38950 19258 38958 19266 sw
rect 70802 19260 71000 19318
tri 38682 19250 38690 19258 ne
rect 38690 19250 38958 19258
tri 38958 19250 38966 19258 sw
tri 38690 19242 38698 19250 ne
rect 38698 19242 38966 19250
tri 38966 19242 38974 19250 sw
tri 38698 19234 38706 19242 ne
rect 38706 19234 38974 19242
tri 38974 19234 38982 19242 sw
tri 38706 19226 38714 19234 ne
rect 38714 19226 38982 19234
tri 38982 19226 38990 19234 sw
tri 38714 19218 38722 19226 ne
rect 38722 19218 38990 19226
tri 38990 19218 38998 19226 sw
tri 38722 19210 38730 19218 ne
rect 38730 19216 38998 19218
rect 38730 19210 38862 19216
tri 38730 19202 38738 19210 ne
rect 38738 19202 38862 19210
tri 38738 19194 38746 19202 ne
rect 38746 19194 38862 19202
tri 38746 19186 38754 19194 ne
rect 38754 19186 38862 19194
tri 38754 19178 38762 19186 ne
rect 38762 19178 38862 19186
tri 38762 19170 38770 19178 ne
rect 38770 19170 38862 19178
rect 38908 19210 38998 19216
tri 38998 19210 39006 19218 sw
rect 70802 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19202 39006 19210
tri 39006 19202 39014 19210 sw
rect 38908 19194 39014 19202
tri 39014 19194 39022 19202 sw
rect 38908 19186 39022 19194
tri 39022 19186 39030 19194 sw
rect 38908 19180 39030 19186
tri 39030 19180 39036 19186 sw
rect 38908 19172 39036 19180
tri 39036 19172 39044 19180 sw
rect 38908 19170 39044 19172
tri 38770 19162 38778 19170 ne
rect 38778 19164 39044 19170
tri 39044 19164 39052 19172 sw
rect 38778 19162 39052 19164
tri 38778 19154 38786 19162 ne
rect 38786 19156 39052 19162
tri 39052 19156 39060 19164 sw
rect 70802 19156 71000 19214
rect 38786 19154 39060 19156
tri 38786 19147 38793 19154 ne
rect 38793 19148 39060 19154
tri 39060 19148 39068 19156 sw
rect 38793 19147 39068 19148
tri 38793 19139 38801 19147 ne
rect 38801 19140 39068 19147
tri 39068 19140 39076 19148 sw
rect 38801 19139 39076 19140
tri 38801 19131 38809 19139 ne
rect 38809 19132 39076 19139
tri 39076 19132 39084 19140 sw
rect 38809 19131 39084 19132
tri 38809 19123 38817 19131 ne
rect 38817 19124 39084 19131
tri 39084 19124 39092 19132 sw
rect 38817 19123 39092 19124
tri 38817 19115 38825 19123 ne
rect 38825 19116 39092 19123
tri 39092 19116 39100 19124 sw
rect 38825 19115 39100 19116
tri 38825 19107 38833 19115 ne
rect 38833 19108 39100 19115
tri 39100 19108 39108 19116 sw
rect 70802 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 38833 19107 39108 19108
tri 39108 19107 39109 19108 sw
tri 38833 19099 38841 19107 ne
rect 38841 19099 39109 19107
tri 39109 19099 39117 19107 sw
tri 38841 19097 38843 19099 ne
rect 38843 19097 39117 19099
tri 38843 19091 38849 19097 ne
rect 38849 19091 39117 19097
tri 39117 19091 39125 19099 sw
tri 38849 19083 38857 19091 ne
rect 38857 19084 39125 19091
rect 38857 19083 38994 19084
tri 38857 19079 38861 19083 ne
rect 38861 19079 38994 19083
tri 38861 19071 38869 19079 ne
rect 38869 19071 38994 19079
tri 38869 19063 38877 19071 ne
rect 38877 19063 38994 19071
tri 38877 19055 38885 19063 ne
rect 38885 19055 38994 19063
tri 38885 19047 38893 19055 ne
rect 38893 19047 38994 19055
tri 38893 19039 38901 19047 ne
rect 38901 19039 38994 19047
tri 38901 19031 38909 19039 ne
rect 38909 19038 38994 19039
rect 39040 19083 39125 19084
tri 39125 19083 39133 19091 sw
rect 39040 19075 39133 19083
tri 39133 19075 39141 19083 sw
rect 39040 19067 39141 19075
tri 39141 19067 39149 19075 sw
rect 39040 19059 39149 19067
tri 39149 19059 39157 19067 sw
rect 39040 19051 39157 19059
tri 39157 19051 39165 19059 sw
rect 70802 19052 71000 19110
rect 39040 19043 39165 19051
tri 39165 19043 39173 19051 sw
rect 39040 19038 39173 19043
rect 38909 19035 39173 19038
tri 39173 19035 39181 19043 sw
rect 38909 19031 39181 19035
tri 38909 19023 38917 19031 ne
rect 38917 19027 39181 19031
tri 39181 19027 39189 19035 sw
rect 38917 19023 39189 19027
tri 38917 19015 38925 19023 ne
rect 38925 19022 39189 19023
tri 39189 19022 39194 19027 sw
rect 38925 19015 39194 19022
tri 38925 19010 38930 19015 ne
rect 38930 19014 39194 19015
tri 39194 19014 39202 19022 sw
rect 38930 19010 39202 19014
tri 38930 19002 38938 19010 ne
rect 38938 19006 39202 19010
tri 39202 19006 39210 19014 sw
rect 70802 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 38938 19002 39210 19006
tri 38938 18994 38946 19002 ne
rect 38946 18998 39210 19002
tri 39210 18998 39218 19006 sw
rect 38946 18994 39218 18998
tri 38946 18986 38954 18994 ne
rect 38954 18990 39218 18994
tri 39218 18990 39226 18998 sw
rect 38954 18986 39226 18990
tri 38954 18978 38962 18986 ne
rect 38962 18982 39226 18986
tri 39226 18982 39234 18990 sw
rect 38962 18978 39234 18982
tri 38962 18970 38970 18978 ne
rect 38970 18974 39234 18978
tri 39234 18974 39242 18982 sw
rect 38970 18970 39242 18974
tri 38970 18962 38978 18970 ne
rect 38978 18966 39242 18970
tri 39242 18966 39250 18974 sw
rect 38978 18962 39250 18966
tri 38978 18954 38986 18962 ne
rect 38986 18958 39250 18962
tri 39250 18958 39258 18966 sw
rect 38986 18954 39258 18958
tri 38986 18946 38994 18954 ne
rect 38994 18952 39258 18954
rect 38994 18946 39126 18952
tri 38994 18938 39002 18946 ne
rect 39002 18938 39126 18946
tri 39002 18930 39010 18938 ne
rect 39010 18930 39126 18938
tri 39010 18922 39018 18930 ne
rect 39018 18922 39126 18930
tri 39018 18914 39026 18922 ne
rect 39026 18914 39126 18922
tri 39026 18906 39034 18914 ne
rect 39034 18906 39126 18914
rect 39172 18950 39258 18952
tri 39258 18950 39266 18958 sw
rect 39172 18942 39266 18950
tri 39266 18942 39274 18950 sw
rect 70802 18948 71000 19006
rect 39172 18934 39274 18942
tri 39274 18934 39282 18942 sw
rect 39172 18926 39282 18934
tri 39282 18926 39290 18934 sw
rect 39172 18918 39290 18926
tri 39290 18918 39298 18926 sw
rect 39172 18910 39298 18918
tri 39298 18910 39306 18918 sw
rect 39172 18906 39306 18910
tri 39034 18898 39042 18906 ne
rect 39042 18902 39306 18906
tri 39306 18902 39314 18910 sw
rect 70802 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
rect 39042 18899 39314 18902
tri 39314 18899 39317 18902 sw
rect 39042 18898 39317 18899
tri 39042 18891 39049 18898 ne
rect 39049 18891 39317 18898
tri 39317 18891 39325 18899 sw
tri 39049 18883 39057 18891 ne
rect 39057 18883 39325 18891
tri 39325 18883 39333 18891 sw
tri 39057 18875 39065 18883 ne
rect 39065 18875 39333 18883
tri 39333 18875 39341 18883 sw
tri 39065 18867 39073 18875 ne
rect 39073 18867 39341 18875
tri 39341 18867 39349 18875 sw
tri 39073 18859 39081 18867 ne
rect 39081 18859 39349 18867
tri 39349 18859 39357 18867 sw
tri 39081 18851 39089 18859 ne
rect 39089 18851 39357 18859
tri 39357 18851 39365 18859 sw
tri 39089 18843 39097 18851 ne
rect 39097 18843 39365 18851
tri 39365 18843 39373 18851 sw
rect 70802 18844 71000 18902
tri 39097 18835 39105 18843 ne
rect 39105 18835 39373 18843
tri 39373 18835 39381 18843 sw
tri 39105 18827 39113 18835 ne
rect 39113 18827 39381 18835
tri 39381 18827 39389 18835 sw
tri 39113 18819 39121 18827 ne
rect 39121 18820 39389 18827
rect 39121 18819 39258 18820
tri 39121 18811 39129 18819 ne
rect 39129 18811 39258 18819
tri 39129 18803 39137 18811 ne
rect 39137 18803 39258 18811
tri 39137 18795 39145 18803 ne
rect 39145 18795 39258 18803
tri 39145 18787 39153 18795 ne
rect 39153 18787 39258 18795
tri 39153 18779 39161 18787 ne
rect 39161 18779 39258 18787
tri 39161 18771 39169 18779 ne
rect 39169 18774 39258 18779
rect 39304 18819 39389 18820
tri 39389 18819 39397 18827 sw
rect 39304 18811 39397 18819
tri 39397 18811 39405 18819 sw
rect 39304 18803 39405 18811
tri 39405 18803 39413 18811 sw
rect 39304 18795 39413 18803
tri 39413 18795 39421 18803 sw
rect 70802 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18787 39421 18795
tri 39421 18787 39429 18795 sw
rect 39304 18779 39429 18787
tri 39429 18779 39437 18787 sw
rect 39304 18774 39437 18779
rect 39169 18771 39437 18774
tri 39437 18771 39445 18779 sw
tri 39169 18763 39177 18771 ne
rect 39177 18763 39445 18771
tri 39445 18763 39453 18771 sw
tri 39177 18762 39178 18763 ne
rect 39178 18762 39453 18763
tri 39178 18754 39186 18762 ne
rect 39186 18755 39453 18762
tri 39453 18755 39461 18763 sw
rect 39186 18754 39461 18755
tri 39186 18746 39194 18754 ne
rect 39194 18747 39461 18754
tri 39461 18747 39469 18755 sw
rect 39194 18746 39469 18747
tri 39194 18738 39202 18746 ne
rect 39202 18739 39469 18746
tri 39469 18739 39477 18747 sw
rect 70802 18740 71000 18798
rect 39202 18738 39477 18739
tri 39202 18730 39210 18738 ne
rect 39210 18731 39477 18738
tri 39477 18731 39485 18739 sw
rect 39210 18730 39485 18731
tri 39210 18722 39218 18730 ne
rect 39218 18723 39485 18730
tri 39485 18723 39493 18731 sw
rect 39218 18722 39493 18723
tri 39218 18714 39226 18722 ne
rect 39226 18715 39493 18722
tri 39493 18715 39501 18723 sw
rect 39226 18714 39501 18715
tri 39226 18706 39234 18714 ne
rect 39234 18707 39501 18714
tri 39501 18707 39509 18715 sw
rect 39234 18706 39509 18707
tri 39234 18698 39242 18706 ne
rect 39242 18699 39509 18706
tri 39509 18699 39517 18707 sw
rect 39242 18698 39517 18699
tri 39242 18690 39250 18698 ne
rect 39250 18691 39517 18698
tri 39517 18691 39525 18699 sw
rect 70802 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 39250 18690 39525 18691
tri 39250 18682 39258 18690 ne
rect 39258 18688 39525 18690
rect 39258 18682 39390 18688
tri 39258 18674 39266 18682 ne
rect 39266 18674 39390 18682
tri 39266 18666 39274 18674 ne
rect 39274 18666 39390 18674
tri 39274 18658 39282 18666 ne
rect 39282 18658 39390 18666
tri 39282 18650 39290 18658 ne
rect 39290 18650 39390 18658
tri 39290 18642 39298 18650 ne
rect 39298 18642 39390 18650
rect 39436 18683 39525 18688
tri 39525 18683 39533 18691 sw
rect 39436 18675 39533 18683
tri 39533 18675 39541 18683 sw
rect 39436 18667 39541 18675
tri 39541 18667 39549 18675 sw
rect 39436 18659 39549 18667
tri 39549 18659 39557 18667 sw
rect 39436 18656 39557 18659
tri 39557 18656 39560 18659 sw
rect 39436 18648 39560 18656
tri 39560 18648 39568 18656 sw
rect 39436 18642 39568 18648
tri 39298 18634 39306 18642 ne
rect 39306 18640 39568 18642
tri 39568 18640 39576 18648 sw
rect 39306 18634 39576 18640
tri 39306 18626 39314 18634 ne
rect 39314 18632 39576 18634
tri 39576 18632 39584 18640 sw
rect 70802 18636 71000 18694
rect 39314 18626 39584 18632
tri 39314 18623 39317 18626 ne
rect 39317 18624 39584 18626
tri 39584 18624 39592 18632 sw
rect 39317 18623 39592 18624
tri 39317 18615 39325 18623 ne
rect 39325 18616 39592 18623
tri 39592 18616 39600 18624 sw
rect 39325 18615 39600 18616
tri 39325 18607 39333 18615 ne
rect 39333 18608 39600 18615
tri 39600 18608 39608 18616 sw
rect 39333 18607 39608 18608
tri 39333 18599 39341 18607 ne
rect 39341 18600 39608 18607
tri 39608 18600 39616 18608 sw
rect 39341 18599 39616 18600
tri 39341 18591 39349 18599 ne
rect 39349 18592 39616 18599
tri 39616 18592 39624 18600 sw
rect 39349 18591 39624 18592
tri 39349 18583 39357 18591 ne
rect 39357 18584 39624 18591
tri 39624 18584 39632 18592 sw
rect 70802 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39357 18583 39632 18584
tri 39357 18575 39365 18583 ne
rect 39365 18576 39632 18583
tri 39632 18576 39640 18584 sw
rect 39365 18575 39640 18576
tri 39640 18575 39641 18576 sw
tri 39365 18567 39373 18575 ne
rect 39373 18567 39641 18575
tri 39641 18567 39649 18575 sw
tri 39373 18559 39381 18567 ne
rect 39381 18559 39649 18567
tri 39649 18559 39657 18567 sw
tri 39381 18555 39385 18559 ne
rect 39385 18556 39657 18559
rect 39385 18555 39522 18556
tri 39385 18551 39389 18555 ne
rect 39389 18551 39522 18555
tri 39389 18543 39397 18551 ne
rect 39397 18543 39522 18551
tri 39397 18535 39405 18543 ne
rect 39405 18535 39522 18543
tri 39405 18527 39413 18535 ne
rect 39413 18527 39522 18535
tri 39413 18519 39421 18527 ne
rect 39421 18519 39522 18527
tri 39421 18511 39429 18519 ne
rect 39429 18511 39522 18519
tri 39429 18503 39437 18511 ne
rect 39437 18510 39522 18511
rect 39568 18551 39657 18556
tri 39657 18551 39665 18559 sw
rect 39568 18543 39665 18551
tri 39665 18543 39673 18551 sw
rect 39568 18535 39673 18543
tri 39673 18535 39681 18543 sw
rect 39568 18527 39681 18535
tri 39681 18527 39689 18535 sw
rect 70802 18532 71000 18590
rect 39568 18519 39689 18527
tri 39689 18519 39697 18527 sw
rect 39568 18511 39697 18519
tri 39697 18511 39705 18519 sw
rect 39568 18510 39705 18511
rect 39437 18503 39705 18510
tri 39705 18503 39713 18511 sw
tri 39437 18495 39445 18503 ne
rect 39445 18495 39713 18503
tri 39713 18495 39721 18503 sw
tri 39445 18487 39453 18495 ne
rect 39453 18487 39721 18495
tri 39721 18487 39729 18495 sw
tri 39453 18482 39458 18487 ne
rect 39458 18482 39729 18487
tri 39458 18474 39466 18482 ne
rect 39466 18479 39729 18482
tri 39729 18479 39737 18487 sw
rect 70802 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39466 18474 39737 18479
tri 39466 18466 39474 18474 ne
rect 39474 18471 39737 18474
tri 39737 18471 39745 18479 sw
rect 39474 18466 39745 18471
tri 39474 18458 39482 18466 ne
rect 39482 18463 39745 18466
tri 39745 18463 39753 18471 sw
rect 39482 18458 39753 18463
tri 39482 18450 39490 18458 ne
rect 39490 18455 39753 18458
tri 39753 18455 39761 18463 sw
rect 39490 18450 39761 18455
tri 39490 18442 39498 18450 ne
rect 39498 18447 39761 18450
tri 39761 18447 39769 18455 sw
rect 39498 18442 39769 18447
tri 39498 18434 39506 18442 ne
rect 39506 18439 39769 18442
tri 39769 18439 39777 18447 sw
rect 39506 18434 39777 18439
tri 39506 18426 39514 18434 ne
rect 39514 18431 39777 18434
tri 39777 18431 39785 18439 sw
rect 39514 18426 39785 18431
tri 39514 18418 39522 18426 ne
rect 39522 18424 39785 18426
rect 39522 18418 39654 18424
tri 39522 18410 39530 18418 ne
rect 39530 18410 39654 18418
tri 39530 18402 39538 18410 ne
rect 39538 18402 39654 18410
tri 39538 18394 39546 18402 ne
rect 39546 18394 39654 18402
tri 39546 18386 39554 18394 ne
rect 39554 18386 39654 18394
tri 39554 18378 39562 18386 ne
rect 39562 18378 39654 18386
rect 39700 18423 39785 18424
tri 39785 18423 39793 18431 sw
rect 70802 18428 71000 18486
rect 39700 18415 39793 18423
tri 39793 18415 39801 18423 sw
rect 39700 18407 39801 18415
tri 39801 18407 39809 18415 sw
rect 39700 18399 39809 18407
tri 39809 18399 39817 18407 sw
rect 39700 18391 39817 18399
tri 39817 18391 39825 18399 sw
rect 39700 18383 39825 18391
tri 39825 18383 39833 18391 sw
rect 39700 18378 39833 18383
tri 39562 18370 39570 18378 ne
rect 39570 18375 39833 18378
tri 39833 18375 39841 18383 sw
rect 70802 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 39570 18370 39841 18375
tri 39570 18362 39578 18370 ne
rect 39578 18367 39841 18370
tri 39841 18367 39849 18375 sw
rect 39578 18362 39849 18367
tri 39578 18354 39586 18362 ne
rect 39586 18360 39849 18362
tri 39849 18360 39856 18367 sw
rect 39586 18354 39856 18360
tri 39586 18352 39588 18354 ne
rect 39588 18352 39856 18354
tri 39856 18352 39864 18360 sw
tri 39588 18344 39596 18352 ne
rect 39596 18344 39864 18352
tri 39864 18344 39872 18352 sw
tri 39596 18336 39604 18344 ne
rect 39604 18336 39872 18344
tri 39872 18336 39880 18344 sw
tri 39604 18328 39612 18336 ne
rect 39612 18328 39880 18336
tri 39880 18328 39888 18336 sw
tri 39612 18320 39620 18328 ne
rect 39620 18320 39888 18328
tri 39888 18320 39896 18328 sw
rect 70802 18324 71000 18382
tri 39620 18312 39628 18320 ne
rect 39628 18312 39896 18320
tri 39896 18312 39904 18320 sw
tri 39628 18304 39636 18312 ne
rect 39636 18304 39904 18312
tri 39904 18304 39912 18312 sw
tri 39636 18296 39644 18304 ne
rect 39644 18296 39912 18304
tri 39912 18296 39920 18304 sw
tri 39644 18288 39652 18296 ne
rect 39652 18292 39920 18296
rect 39652 18288 39786 18292
tri 39652 18280 39660 18288 ne
rect 39660 18280 39786 18288
tri 39660 18275 39665 18280 ne
rect 39665 18275 39786 18280
tri 39665 18267 39673 18275 ne
rect 39673 18267 39786 18275
tri 39673 18259 39681 18267 ne
rect 39681 18259 39786 18267
tri 39681 18251 39689 18259 ne
rect 39689 18251 39786 18259
tri 39689 18243 39697 18251 ne
rect 39697 18246 39786 18251
rect 39832 18288 39920 18292
tri 39920 18288 39928 18296 sw
rect 39832 18280 39928 18288
tri 39928 18280 39936 18288 sw
rect 39832 18275 39936 18280
tri 39936 18275 39941 18280 sw
rect 70802 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 39832 18267 39941 18275
tri 39941 18267 39949 18275 sw
rect 39832 18259 39949 18267
tri 39949 18259 39957 18267 sw
rect 39832 18251 39957 18259
tri 39957 18251 39965 18259 sw
rect 39832 18246 39965 18251
rect 39697 18243 39965 18246
tri 39965 18243 39973 18251 sw
tri 39697 18235 39705 18243 ne
rect 39705 18235 39973 18243
tri 39973 18235 39981 18243 sw
tri 39705 18227 39713 18235 ne
rect 39713 18227 39981 18235
tri 39981 18227 39989 18235 sw
tri 39713 18219 39721 18227 ne
rect 39721 18219 39989 18227
tri 39989 18219 39997 18227 sw
rect 70802 18220 71000 18278
tri 39721 18211 39729 18219 ne
rect 39729 18211 39997 18219
tri 39997 18211 40005 18219 sw
tri 39729 18203 39737 18211 ne
rect 39737 18203 40005 18211
tri 40005 18203 40013 18211 sw
tri 39737 18195 39745 18203 ne
rect 39745 18195 40013 18203
tri 40013 18195 40021 18203 sw
tri 39745 18187 39753 18195 ne
rect 39753 18187 40021 18195
tri 40021 18187 40029 18195 sw
tri 39753 18179 39761 18187 ne
rect 39761 18179 40029 18187
tri 40029 18179 40037 18187 sw
tri 39761 18171 39769 18179 ne
rect 39769 18171 40037 18179
tri 40037 18171 40045 18179 sw
rect 70802 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
tri 39769 18163 39777 18171 ne
rect 39777 18163 40045 18171
tri 40045 18163 40053 18171 sw
tri 39777 18161 39779 18163 ne
rect 39779 18161 40053 18163
tri 40053 18161 40055 18163 sw
tri 39779 18153 39787 18161 ne
rect 39787 18160 40055 18161
rect 39787 18153 39918 18160
tri 39787 18145 39795 18153 ne
rect 39795 18145 39918 18153
tri 39795 18137 39803 18145 ne
rect 39803 18137 39918 18145
tri 39803 18129 39811 18137 ne
rect 39811 18129 39918 18137
tri 39811 18121 39819 18129 ne
rect 39819 18121 39918 18129
tri 39819 18113 39827 18121 ne
rect 39827 18114 39918 18121
rect 39964 18153 40055 18160
tri 40055 18153 40063 18161 sw
rect 39964 18145 40063 18153
tri 40063 18145 40071 18153 sw
rect 39964 18137 40071 18145
tri 40071 18137 40079 18145 sw
rect 39964 18129 40079 18137
tri 40079 18129 40087 18137 sw
rect 39964 18121 40087 18129
tri 40087 18121 40095 18129 sw
rect 39964 18114 40095 18121
rect 39827 18113 40095 18114
tri 40095 18113 40103 18121 sw
rect 70802 18116 71000 18174
tri 39827 18105 39835 18113 ne
rect 39835 18105 40103 18113
tri 40103 18105 40111 18113 sw
tri 39835 18097 39843 18105 ne
rect 39843 18097 40111 18105
tri 40111 18097 40119 18105 sw
tri 39843 18089 39851 18097 ne
rect 39851 18089 40119 18097
tri 40119 18089 40127 18097 sw
tri 39851 18081 39859 18089 ne
rect 39859 18081 40127 18089
tri 40127 18081 40135 18089 sw
tri 39859 18073 39867 18081 ne
rect 39867 18073 40135 18081
tri 40135 18073 40143 18081 sw
tri 39867 18065 39875 18073 ne
rect 39875 18065 40143 18073
tri 40143 18065 40151 18073 sw
rect 70802 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39875 18057 39883 18065 ne
rect 39883 18057 40151 18065
tri 40151 18057 40159 18065 sw
tri 39883 18049 39891 18057 ne
rect 39891 18049 40159 18057
tri 40159 18049 40167 18057 sw
tri 39891 18047 39893 18049 ne
rect 39893 18047 40167 18049
tri 40167 18047 40169 18049 sw
tri 39893 18039 39901 18047 ne
rect 39901 18039 40169 18047
tri 40169 18039 40177 18047 sw
tri 39901 18031 39909 18039 ne
rect 39909 18031 40177 18039
tri 40177 18031 40185 18039 sw
tri 39909 18023 39917 18031 ne
rect 39917 18028 40185 18031
rect 39917 18023 40050 18028
tri 39917 18015 39925 18023 ne
rect 39925 18015 40050 18023
tri 39925 18007 39933 18015 ne
rect 39933 18007 40050 18015
tri 39933 17999 39941 18007 ne
rect 39941 17999 40050 18007
tri 39941 17991 39949 17999 ne
rect 39949 17991 40050 17999
tri 39949 17983 39957 17991 ne
rect 39957 17983 40050 17991
tri 39957 17975 39965 17983 ne
rect 39965 17982 40050 17983
rect 40096 18023 40185 18028
tri 40185 18023 40193 18031 sw
rect 40096 18015 40193 18023
tri 40193 18015 40201 18023 sw
rect 40096 18007 40201 18015
tri 40201 18007 40209 18015 sw
rect 70802 18012 71000 18070
rect 40096 17999 40209 18007
tri 40209 17999 40217 18007 sw
rect 40096 17991 40217 17999
tri 40217 17991 40225 17999 sw
rect 40096 17983 40225 17991
tri 40225 17983 40233 17991 sw
rect 40096 17982 40233 17983
rect 39965 17975 40233 17982
tri 40233 17975 40241 17983 sw
tri 39965 17967 39973 17975 ne
rect 39973 17969 40241 17975
tri 40241 17969 40247 17975 sw
rect 39973 17967 40247 17969
tri 39973 17959 39981 17967 ne
rect 39981 17961 40247 17967
tri 40247 17961 40255 17969 sw
rect 70802 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 39981 17959 40255 17961
tri 39981 17951 39989 17959 ne
rect 39989 17953 40255 17959
tri 40255 17953 40263 17961 sw
rect 39989 17951 40263 17953
tri 39989 17943 39997 17951 ne
rect 39997 17945 40263 17951
tri 40263 17945 40271 17953 sw
rect 39997 17943 40271 17945
tri 39997 17935 40005 17943 ne
rect 40005 17937 40271 17943
tri 40271 17937 40279 17945 sw
rect 40005 17935 40279 17937
tri 40005 17927 40013 17935 ne
rect 40013 17929 40279 17935
tri 40279 17929 40287 17937 sw
rect 40013 17927 40287 17929
tri 40013 17919 40021 17927 ne
rect 40021 17921 40287 17927
tri 40287 17921 40295 17929 sw
rect 40021 17919 40295 17921
tri 40021 17911 40029 17919 ne
rect 40029 17913 40295 17919
tri 40295 17913 40303 17921 sw
rect 40029 17911 40303 17913
tri 40029 17909 40031 17911 ne
rect 40031 17909 40303 17911
tri 40031 17901 40039 17909 ne
rect 40039 17905 40303 17909
tri 40303 17905 40311 17913 sw
rect 70802 17908 71000 17966
rect 40039 17901 40311 17905
tri 40039 17893 40047 17901 ne
rect 40047 17897 40311 17901
tri 40311 17897 40319 17905 sw
rect 40047 17896 40319 17897
rect 40047 17893 40182 17896
tri 40047 17885 40055 17893 ne
rect 40055 17885 40182 17893
tri 40055 17877 40063 17885 ne
rect 40063 17877 40182 17885
tri 40063 17869 40071 17877 ne
rect 40071 17869 40182 17877
tri 40071 17861 40079 17869 ne
rect 40079 17861 40182 17869
tri 40079 17853 40087 17861 ne
rect 40087 17853 40182 17861
tri 40087 17845 40095 17853 ne
rect 40095 17850 40182 17853
rect 40228 17889 40319 17896
tri 40319 17889 40327 17897 sw
rect 40228 17881 40327 17889
tri 40327 17881 40335 17889 sw
rect 40228 17873 40335 17881
tri 40335 17873 40343 17881 sw
rect 40228 17865 40343 17873
tri 40343 17865 40351 17873 sw
rect 40228 17857 40351 17865
tri 40351 17857 40359 17865 sw
rect 70802 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 40228 17850 40359 17857
rect 40095 17849 40359 17850
tri 40359 17849 40367 17857 sw
rect 40095 17845 40367 17849
tri 40095 17837 40103 17845 ne
rect 40103 17841 40367 17845
tri 40367 17841 40375 17849 sw
rect 40103 17837 40375 17841
tri 40103 17829 40111 17837 ne
rect 40111 17833 40375 17837
tri 40375 17833 40383 17841 sw
rect 40111 17829 40383 17833
tri 40111 17821 40119 17829 ne
rect 40119 17827 40383 17829
tri 40383 17827 40389 17833 sw
rect 40119 17821 40389 17827
tri 40119 17813 40127 17821 ne
rect 40127 17819 40389 17821
tri 40389 17819 40397 17827 sw
rect 40127 17813 40397 17819
tri 40127 17805 40135 17813 ne
rect 40135 17811 40397 17813
tri 40397 17811 40405 17819 sw
rect 40135 17805 40405 17811
tri 40135 17797 40143 17805 ne
rect 40143 17803 40405 17805
tri 40405 17803 40413 17811 sw
rect 70802 17804 71000 17862
rect 40143 17797 40413 17803
tri 40143 17789 40151 17797 ne
rect 40151 17795 40413 17797
tri 40413 17795 40421 17803 sw
rect 40151 17789 40421 17795
tri 40151 17781 40159 17789 ne
rect 40159 17787 40421 17789
tri 40421 17787 40429 17795 sw
rect 40159 17781 40429 17787
tri 40159 17773 40167 17781 ne
rect 40167 17779 40429 17781
tri 40429 17779 40437 17787 sw
rect 40167 17773 40437 17779
tri 40167 17765 40175 17773 ne
rect 40175 17771 40437 17773
tri 40437 17771 40445 17779 sw
rect 40175 17765 40445 17771
tri 40175 17763 40177 17765 ne
rect 40177 17764 40445 17765
rect 40177 17763 40314 17764
tri 40177 17755 40185 17763 ne
rect 40185 17755 40314 17763
tri 40185 17747 40193 17755 ne
rect 40193 17747 40314 17755
tri 40193 17739 40201 17747 ne
rect 40201 17739 40314 17747
tri 40201 17731 40209 17739 ne
rect 40209 17731 40314 17739
tri 40209 17723 40217 17731 ne
rect 40217 17723 40314 17731
tri 40217 17715 40225 17723 ne
rect 40225 17718 40314 17723
rect 40360 17763 40445 17764
tri 40445 17763 40453 17771 sw
rect 40360 17755 40453 17763
tri 40453 17755 40461 17763 sw
rect 70802 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17747 40461 17755
tri 40461 17747 40469 17755 sw
rect 40360 17739 40469 17747
tri 40469 17739 40477 17747 sw
rect 40360 17731 40477 17739
tri 40477 17731 40485 17739 sw
rect 40360 17723 40485 17731
tri 40485 17723 40493 17731 sw
rect 40360 17718 40493 17723
rect 40225 17715 40493 17718
tri 40493 17715 40501 17723 sw
tri 40225 17707 40233 17715 ne
rect 40233 17707 40501 17715
tri 40501 17707 40509 17715 sw
tri 40233 17699 40241 17707 ne
rect 40241 17699 40509 17707
tri 40509 17699 40517 17707 sw
rect 70802 17700 71000 17758
tri 40241 17691 40249 17699 ne
rect 40249 17691 40517 17699
tri 40517 17691 40525 17699 sw
tri 40249 17685 40255 17691 ne
rect 40255 17688 40525 17691
tri 40525 17688 40528 17691 sw
rect 40255 17685 40528 17688
tri 40255 17677 40263 17685 ne
rect 40263 17680 40528 17685
tri 40528 17680 40536 17688 sw
rect 40263 17677 40536 17680
tri 40263 17669 40271 17677 ne
rect 40271 17672 40536 17677
tri 40536 17672 40544 17680 sw
rect 40271 17669 40544 17672
tri 40271 17661 40279 17669 ne
rect 40279 17664 40544 17669
tri 40544 17664 40552 17672 sw
rect 40279 17661 40552 17664
tri 40279 17653 40287 17661 ne
rect 40287 17656 40552 17661
tri 40552 17656 40560 17664 sw
rect 40287 17653 40560 17656
tri 40287 17645 40295 17653 ne
rect 40295 17648 40560 17653
tri 40560 17648 40568 17656 sw
rect 70802 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
rect 40295 17645 40568 17648
tri 40295 17637 40303 17645 ne
rect 40303 17640 40568 17645
tri 40568 17640 40576 17648 sw
rect 40303 17637 40576 17640
tri 40303 17629 40311 17637 ne
rect 40311 17632 40576 17637
tri 40576 17632 40584 17640 sw
rect 40311 17629 40446 17632
tri 40311 17621 40319 17629 ne
rect 40319 17621 40446 17629
tri 40319 17613 40327 17621 ne
rect 40327 17613 40446 17621
tri 40327 17605 40335 17613 ne
rect 40335 17605 40446 17613
tri 40335 17597 40343 17605 ne
rect 40343 17597 40446 17605
tri 40343 17589 40351 17597 ne
rect 40351 17589 40446 17597
tri 40351 17581 40359 17589 ne
rect 40359 17586 40446 17589
rect 40492 17624 40584 17632
tri 40584 17624 40592 17632 sw
rect 40492 17616 40592 17624
tri 40592 17616 40600 17624 sw
rect 40492 17608 40600 17616
tri 40600 17608 40608 17616 sw
rect 40492 17600 40608 17608
tri 40608 17600 40616 17608 sw
rect 40492 17592 40616 17600
tri 40616 17592 40624 17600 sw
rect 70802 17596 71000 17654
rect 40492 17586 40624 17592
rect 40359 17584 40624 17586
tri 40624 17584 40632 17592 sw
rect 40359 17581 40632 17584
tri 40359 17573 40367 17581 ne
rect 40367 17578 40632 17581
tri 40632 17578 40638 17584 sw
rect 40367 17573 40638 17578
tri 40367 17570 40370 17573 ne
rect 40370 17570 40638 17573
tri 40638 17570 40646 17578 sw
tri 40370 17562 40378 17570 ne
rect 40378 17562 40646 17570
tri 40646 17562 40654 17570 sw
tri 40378 17554 40386 17562 ne
rect 40386 17554 40654 17562
tri 40654 17554 40662 17562 sw
tri 40386 17546 40394 17554 ne
rect 40394 17546 40662 17554
tri 40662 17546 40670 17554 sw
rect 70802 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
tri 40394 17538 40402 17546 ne
rect 40402 17538 40670 17546
tri 40670 17538 40678 17546 sw
tri 40402 17530 40410 17538 ne
rect 40410 17530 40678 17538
tri 40678 17530 40686 17538 sw
tri 40410 17522 40418 17530 ne
rect 40418 17522 40686 17530
tri 40686 17522 40694 17530 sw
tri 40418 17514 40426 17522 ne
rect 40426 17514 40694 17522
tri 40694 17514 40702 17522 sw
tri 40426 17506 40434 17514 ne
rect 40434 17506 40702 17514
tri 40702 17506 40710 17514 sw
tri 40434 17502 40438 17506 ne
rect 40438 17502 40710 17506
tri 40710 17502 40714 17506 sw
tri 40438 17498 40442 17502 ne
rect 40442 17500 40714 17502
rect 40442 17498 40578 17500
tri 40442 17490 40450 17498 ne
rect 40450 17490 40578 17498
tri 40450 17482 40458 17490 ne
rect 40458 17482 40578 17490
tri 40458 17474 40466 17482 ne
rect 40466 17474 40578 17482
tri 40466 17466 40474 17474 ne
rect 40474 17466 40578 17474
tri 40474 17458 40482 17466 ne
rect 40482 17458 40578 17466
tri 40482 17450 40490 17458 ne
rect 40490 17454 40578 17458
rect 40624 17498 40714 17500
tri 40714 17498 40718 17502 sw
rect 40624 17490 40718 17498
tri 40718 17490 40726 17498 sw
rect 70802 17492 71000 17550
rect 40624 17482 40726 17490
tri 40726 17482 40734 17490 sw
rect 40624 17474 40734 17482
tri 40734 17474 40742 17482 sw
rect 40624 17466 40742 17474
tri 40742 17466 40750 17474 sw
rect 40624 17458 40750 17466
tri 40750 17458 40758 17466 sw
rect 40624 17454 40758 17458
rect 40490 17450 40758 17454
tri 40758 17450 40766 17458 sw
tri 40490 17442 40498 17450 ne
rect 40498 17442 40766 17450
tri 40766 17442 40774 17450 sw
rect 70802 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
tri 40498 17434 40506 17442 ne
rect 40506 17434 40774 17442
tri 40774 17434 40782 17442 sw
tri 40506 17426 40514 17434 ne
rect 40514 17426 40782 17434
tri 40782 17426 40790 17434 sw
tri 40514 17418 40522 17426 ne
rect 40522 17418 40790 17426
tri 40790 17418 40798 17426 sw
tri 40522 17410 40530 17418 ne
rect 40530 17410 40798 17418
tri 40798 17410 40806 17418 sw
tri 40530 17402 40538 17410 ne
rect 40538 17402 40806 17410
tri 40806 17402 40814 17410 sw
tri 40538 17394 40546 17402 ne
rect 40546 17394 40814 17402
tri 40814 17394 40822 17402 sw
tri 40546 17386 40554 17394 ne
rect 40554 17386 40822 17394
tri 40822 17386 40830 17394 sw
rect 70802 17388 71000 17446
tri 40554 17378 40562 17386 ne
rect 40562 17378 40830 17386
tri 40830 17378 40838 17386 sw
tri 40562 17370 40570 17378 ne
rect 40570 17370 40838 17378
tri 40838 17370 40846 17378 sw
tri 40570 17365 40575 17370 ne
rect 40575 17368 40846 17370
rect 40575 17365 40710 17368
tri 40575 17357 40583 17365 ne
rect 40583 17357 40710 17365
tri 40583 17349 40591 17357 ne
rect 40591 17349 40710 17357
tri 40591 17341 40599 17349 ne
rect 40599 17341 40710 17349
tri 40599 17333 40607 17341 ne
rect 40607 17333 40710 17341
tri 40607 17325 40615 17333 ne
rect 40615 17325 40710 17333
tri 40615 17317 40623 17325 ne
rect 40623 17322 40710 17325
rect 40756 17365 40846 17368
tri 40846 17365 40851 17370 sw
rect 40756 17357 40851 17365
tri 40851 17357 40859 17365 sw
rect 40756 17349 40859 17357
tri 40859 17349 40867 17357 sw
rect 40756 17341 40867 17349
tri 40867 17341 40875 17349 sw
rect 70802 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17333 40875 17341
tri 40875 17333 40883 17341 sw
rect 40756 17325 40883 17333
tri 40883 17325 40891 17333 sw
rect 40756 17322 40891 17325
rect 40623 17317 40891 17322
tri 40891 17317 40899 17325 sw
tri 40623 17309 40631 17317 ne
rect 40631 17309 40899 17317
tri 40899 17309 40907 17317 sw
tri 40631 17301 40639 17309 ne
rect 40639 17301 40907 17309
tri 40907 17301 40915 17309 sw
tri 40639 17293 40647 17301 ne
rect 40647 17293 40915 17301
tri 40915 17293 40923 17301 sw
tri 40647 17285 40655 17293 ne
rect 40655 17285 40923 17293
tri 40923 17285 40931 17293 sw
tri 40655 17277 40663 17285 ne
rect 40663 17277 40931 17285
tri 40931 17277 40939 17285 sw
rect 70802 17284 71000 17342
tri 40663 17269 40671 17277 ne
rect 40671 17269 40939 17277
tri 40939 17269 40947 17277 sw
tri 40671 17261 40679 17269 ne
rect 40679 17261 40947 17269
tri 40947 17261 40955 17269 sw
tri 40679 17253 40687 17261 ne
rect 40687 17253 40955 17261
tri 40955 17253 40963 17261 sw
tri 40687 17245 40695 17253 ne
rect 40695 17245 40963 17253
tri 40963 17245 40971 17253 sw
tri 40695 17237 40703 17245 ne
rect 40703 17237 40971 17245
tri 40971 17237 40979 17245 sw
rect 70802 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
tri 40703 17229 40711 17237 ne
rect 40711 17236 40979 17237
rect 40711 17229 40842 17236
tri 40711 17227 40713 17229 ne
rect 40713 17227 40842 17229
tri 40713 17222 40718 17227 ne
rect 40718 17222 40842 17227
tri 40718 17219 40721 17222 ne
rect 40721 17219 40842 17222
tri 40721 17211 40729 17219 ne
rect 40729 17211 40842 17219
tri 40729 17203 40737 17211 ne
rect 40737 17203 40842 17211
tri 40737 17195 40745 17203 ne
rect 40745 17195 40842 17203
tri 40745 17187 40753 17195 ne
rect 40753 17190 40842 17195
rect 40888 17229 40979 17236
tri 40979 17229 40987 17237 sw
rect 40888 17227 40987 17229
tri 40987 17227 40989 17229 sw
rect 40888 17219 40989 17227
tri 40989 17219 40997 17227 sw
rect 40888 17211 40997 17219
tri 40997 17211 41005 17219 sw
rect 40888 17203 41005 17211
tri 41005 17203 41013 17211 sw
rect 40888 17195 41013 17203
tri 41013 17195 41021 17203 sw
rect 40888 17190 41021 17195
rect 40753 17187 41021 17190
tri 41021 17187 41029 17195 sw
tri 40753 17179 40761 17187 ne
rect 40761 17179 41029 17187
tri 41029 17179 41037 17187 sw
rect 70802 17180 71000 17238
tri 40761 17171 40769 17179 ne
rect 40769 17171 41037 17179
tri 41037 17171 41045 17179 sw
tri 40769 17163 40777 17171 ne
rect 40777 17163 41045 17171
tri 41045 17163 41053 17171 sw
tri 40777 17155 40785 17163 ne
rect 40785 17155 41053 17163
tri 41053 17155 41061 17163 sw
tri 40785 17147 40793 17155 ne
rect 40793 17147 41061 17155
tri 41061 17147 41069 17155 sw
tri 40793 17139 40801 17147 ne
rect 40801 17139 41069 17147
tri 41069 17139 41077 17147 sw
tri 40801 17131 40809 17139 ne
rect 40809 17131 41077 17139
tri 41077 17131 41085 17139 sw
rect 70802 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40809 17123 40817 17131 ne
rect 40817 17123 41085 17131
tri 41085 17123 41093 17131 sw
tri 40817 17115 40825 17123 ne
rect 40825 17115 41093 17123
tri 41093 17115 41101 17123 sw
tri 40825 17107 40833 17115 ne
rect 40833 17110 41101 17115
tri 41101 17110 41106 17115 sw
rect 40833 17107 41106 17110
tri 40833 17099 40841 17107 ne
rect 40841 17104 41106 17107
rect 40841 17099 40974 17104
tri 40841 17091 40849 17099 ne
rect 40849 17091 40974 17099
tri 40849 17090 40850 17091 ne
rect 40850 17090 40974 17091
tri 40850 17082 40858 17090 ne
rect 40858 17082 40974 17090
tri 40858 17074 40866 17082 ne
rect 40866 17074 40974 17082
tri 40866 17066 40874 17074 ne
rect 40874 17066 40974 17074
tri 40874 17058 40882 17066 ne
rect 40882 17058 40974 17066
rect 41020 17102 41106 17104
tri 41106 17102 41114 17110 sw
rect 41020 17094 41114 17102
tri 41114 17094 41122 17102 sw
rect 41020 17086 41122 17094
tri 41122 17086 41130 17094 sw
rect 41020 17078 41130 17086
tri 41130 17078 41138 17086 sw
rect 41020 17070 41138 17078
tri 41138 17070 41146 17078 sw
rect 70802 17076 71000 17134
rect 41020 17062 41146 17070
tri 41146 17062 41154 17070 sw
rect 41020 17058 41154 17062
tri 40882 17050 40890 17058 ne
rect 40890 17054 41154 17058
tri 41154 17054 41162 17062 sw
rect 40890 17050 41162 17054
tri 40890 17042 40898 17050 ne
rect 40898 17046 41162 17050
tri 41162 17046 41170 17054 sw
rect 40898 17042 41170 17046
tri 40898 17034 40906 17042 ne
rect 40906 17038 41170 17042
tri 41170 17038 41178 17046 sw
rect 40906 17034 41178 17038
tri 40906 17026 40914 17034 ne
rect 40914 17030 41178 17034
tri 41178 17030 41186 17038 sw
rect 70802 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 40914 17026 41186 17030
tri 40914 17018 40922 17026 ne
rect 40922 17022 41186 17026
tri 41186 17022 41194 17030 sw
rect 40922 17018 41194 17022
tri 40922 17010 40930 17018 ne
rect 40930 17014 41194 17018
tri 41194 17014 41202 17022 sw
rect 40930 17010 41202 17014
tri 40930 17002 40938 17010 ne
rect 40938 17006 41202 17010
tri 41202 17006 41210 17014 sw
rect 40938 17002 41210 17006
tri 40938 16994 40946 17002 ne
rect 40946 16999 41210 17002
tri 41210 16999 41217 17006 sw
rect 40946 16994 41217 16999
tri 40946 16986 40954 16994 ne
rect 40954 16991 41217 16994
tri 41217 16991 41225 16999 sw
rect 40954 16986 41225 16991
tri 40954 16978 40962 16986 ne
rect 40962 16983 41225 16986
tri 41225 16983 41233 16991 sw
rect 40962 16978 41233 16983
tri 40962 16970 40970 16978 ne
rect 40970 16975 41233 16978
tri 41233 16975 41241 16983 sw
rect 40970 16972 41241 16975
rect 40970 16970 41106 16972
tri 40970 16966 40974 16970 ne
rect 40974 16966 41106 16970
tri 40974 16962 40978 16966 ne
rect 40978 16962 41106 16966
tri 40978 16954 40986 16962 ne
rect 40986 16954 41106 16962
tri 40986 16946 40994 16954 ne
rect 40994 16946 41106 16954
tri 40994 16938 41002 16946 ne
rect 41002 16938 41106 16946
tri 41002 16930 41010 16938 ne
rect 41010 16930 41106 16938
tri 41010 16922 41018 16930 ne
rect 41018 16926 41106 16930
rect 41152 16970 41241 16972
tri 41241 16970 41246 16975 sw
rect 70802 16972 71000 17030
rect 41152 16962 41246 16970
tri 41246 16962 41254 16970 sw
rect 41152 16954 41254 16962
tri 41254 16954 41262 16962 sw
rect 41152 16946 41262 16954
tri 41262 16946 41270 16954 sw
rect 41152 16938 41270 16946
tri 41270 16938 41278 16946 sw
rect 41152 16930 41278 16938
tri 41278 16930 41286 16938 sw
rect 41152 16926 41286 16930
rect 41018 16922 41286 16926
tri 41286 16922 41294 16930 sw
rect 70802 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41018 16914 41026 16922 ne
rect 41026 16914 41294 16922
tri 41294 16914 41302 16922 sw
tri 41026 16906 41034 16914 ne
rect 41034 16908 41302 16914
tri 41302 16908 41308 16914 sw
rect 41034 16906 41308 16908
tri 41034 16898 41042 16906 ne
rect 41042 16900 41308 16906
tri 41308 16900 41316 16908 sw
rect 41042 16898 41316 16900
tri 41042 16890 41050 16898 ne
rect 41050 16892 41316 16898
tri 41316 16892 41324 16900 sw
rect 41050 16890 41324 16892
tri 41050 16882 41058 16890 ne
rect 41058 16884 41324 16890
tri 41324 16884 41332 16892 sw
rect 41058 16882 41332 16884
tri 41058 16874 41066 16882 ne
rect 41066 16876 41332 16882
tri 41332 16876 41340 16884 sw
rect 41066 16874 41340 16876
tri 41066 16866 41074 16874 ne
rect 41074 16868 41340 16874
tri 41340 16868 41348 16876 sw
rect 70802 16868 71000 16926
rect 41074 16866 41348 16868
tri 41074 16858 41082 16866 ne
rect 41082 16860 41348 16866
tri 41348 16860 41356 16868 sw
rect 41082 16858 41356 16860
tri 41082 16850 41090 16858 ne
rect 41090 16852 41356 16858
tri 41356 16852 41364 16860 sw
rect 41090 16850 41364 16852
tri 41090 16842 41098 16850 ne
rect 41098 16844 41364 16850
tri 41364 16844 41372 16852 sw
rect 41098 16842 41372 16844
tri 41098 16834 41106 16842 ne
rect 41106 16840 41372 16842
rect 41106 16834 41238 16840
tri 41106 16826 41114 16834 ne
rect 41114 16826 41238 16834
tri 41114 16818 41122 16826 ne
rect 41122 16818 41238 16826
tri 41122 16810 41130 16818 ne
rect 41130 16810 41238 16818
tri 41130 16802 41138 16810 ne
rect 41138 16802 41238 16810
tri 41138 16794 41146 16802 ne
rect 41146 16794 41238 16802
rect 41284 16836 41372 16840
tri 41372 16836 41380 16844 sw
rect 41284 16828 41380 16836
tri 41380 16828 41388 16836 sw
rect 41284 16820 41388 16828
tri 41388 16820 41396 16828 sw
rect 70802 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16812 41396 16820
tri 41396 16812 41404 16820 sw
rect 41284 16804 41404 16812
tri 41404 16804 41412 16812 sw
rect 41284 16796 41412 16804
tri 41412 16796 41420 16804 sw
rect 41284 16794 41420 16796
tri 41146 16786 41154 16794 ne
rect 41154 16789 41420 16794
tri 41420 16789 41427 16796 sw
rect 41154 16786 41427 16789
tri 41154 16778 41162 16786 ne
rect 41162 16781 41427 16786
tri 41427 16781 41435 16789 sw
rect 41162 16778 41435 16781
tri 41162 16770 41170 16778 ne
rect 41170 16773 41435 16778
tri 41435 16773 41443 16781 sw
rect 41170 16770 41443 16773
tri 41170 16763 41177 16770 ne
rect 41177 16765 41443 16770
tri 41443 16765 41451 16773 sw
rect 41177 16763 41451 16765
tri 41177 16755 41185 16763 ne
rect 41185 16757 41451 16763
tri 41451 16757 41459 16765 sw
rect 70802 16764 71000 16822
rect 41185 16755 41459 16757
tri 41185 16747 41193 16755 ne
rect 41193 16749 41459 16755
tri 41459 16749 41467 16757 sw
rect 41193 16747 41467 16749
tri 41193 16739 41201 16747 ne
rect 41201 16741 41467 16747
tri 41467 16741 41475 16749 sw
rect 41201 16739 41475 16741
tri 41201 16731 41209 16739 ne
rect 41209 16733 41475 16739
tri 41475 16733 41483 16741 sw
rect 41209 16731 41483 16733
tri 41209 16723 41217 16731 ne
rect 41217 16725 41483 16731
tri 41483 16725 41491 16733 sw
rect 41217 16723 41491 16725
tri 41217 16715 41225 16723 ne
rect 41225 16717 41491 16723
tri 41491 16717 41499 16725 sw
rect 70802 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 41225 16715 41499 16717
tri 41499 16715 41501 16717 sw
tri 41225 16707 41233 16715 ne
rect 41233 16708 41501 16715
rect 41233 16707 41370 16708
tri 41233 16702 41238 16707 ne
rect 41238 16702 41370 16707
tri 41238 16699 41241 16702 ne
rect 41241 16699 41370 16702
tri 41241 16691 41249 16699 ne
rect 41249 16691 41370 16699
tri 41249 16683 41257 16691 ne
rect 41257 16683 41370 16691
tri 41257 16675 41265 16683 ne
rect 41265 16675 41370 16683
tri 41265 16667 41273 16675 ne
rect 41273 16667 41370 16675
tri 41273 16659 41281 16667 ne
rect 41281 16662 41370 16667
rect 41416 16707 41501 16708
tri 41501 16707 41509 16715 sw
rect 41416 16699 41509 16707
tri 41509 16699 41517 16707 sw
rect 41416 16691 41517 16699
tri 41517 16691 41525 16699 sw
rect 41416 16683 41525 16691
tri 41525 16683 41533 16691 sw
rect 41416 16675 41533 16683
tri 41533 16675 41541 16683 sw
rect 41416 16667 41541 16675
tri 41541 16667 41549 16675 sw
rect 41416 16662 41549 16667
rect 41281 16659 41549 16662
tri 41549 16659 41557 16667 sw
rect 70802 16660 71000 16718
tri 41281 16651 41289 16659 ne
rect 41289 16651 41557 16659
tri 41557 16651 41565 16659 sw
tri 41289 16643 41297 16651 ne
rect 41297 16643 41565 16651
tri 41565 16643 41573 16651 sw
tri 41297 16635 41305 16643 ne
rect 41305 16638 41573 16643
tri 41573 16638 41578 16643 sw
rect 41305 16635 41578 16638
tri 41305 16634 41306 16635 ne
rect 41306 16634 41578 16635
tri 41306 16626 41314 16634 ne
rect 41314 16630 41578 16634
tri 41578 16630 41586 16638 sw
rect 41314 16626 41586 16630
tri 41314 16618 41322 16626 ne
rect 41322 16622 41586 16626
tri 41586 16622 41594 16630 sw
rect 41322 16618 41594 16622
tri 41322 16610 41330 16618 ne
rect 41330 16614 41594 16618
tri 41594 16614 41602 16622 sw
rect 70802 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41330 16610 41602 16614
tri 41330 16602 41338 16610 ne
rect 41338 16606 41602 16610
tri 41602 16606 41610 16614 sw
rect 41338 16602 41610 16606
tri 41338 16594 41346 16602 ne
rect 41346 16598 41610 16602
tri 41610 16598 41618 16606 sw
rect 41346 16594 41618 16598
tri 41346 16586 41354 16594 ne
rect 41354 16590 41618 16594
tri 41618 16590 41626 16598 sw
rect 41354 16586 41626 16590
tri 41354 16578 41362 16586 ne
rect 41362 16582 41626 16586
tri 41626 16582 41634 16590 sw
rect 41362 16578 41634 16582
tri 41362 16570 41370 16578 ne
rect 41370 16576 41634 16578
rect 41370 16570 41502 16576
tri 41370 16562 41378 16570 ne
rect 41378 16562 41502 16570
tri 41378 16554 41386 16562 ne
rect 41386 16554 41502 16562
tri 41386 16546 41394 16554 ne
rect 41394 16546 41502 16554
tri 41394 16538 41402 16546 ne
rect 41402 16538 41502 16546
tri 41402 16530 41410 16538 ne
rect 41410 16530 41502 16538
rect 41548 16574 41634 16576
tri 41634 16574 41642 16582 sw
rect 41548 16566 41642 16574
tri 41642 16566 41650 16574 sw
rect 41548 16558 41650 16566
tri 41650 16558 41658 16566 sw
rect 41548 16550 41658 16558
tri 41658 16550 41666 16558 sw
rect 70802 16556 71000 16614
rect 41548 16542 41666 16550
tri 41666 16542 41674 16550 sw
rect 41548 16534 41674 16542
tri 41674 16534 41682 16542 sw
rect 41548 16530 41682 16534
tri 41410 16522 41418 16530 ne
rect 41418 16526 41682 16530
tri 41682 16526 41690 16534 sw
rect 41418 16522 41690 16526
tri 41690 16522 41694 16526 sw
tri 41418 16514 41426 16522 ne
rect 41426 16514 41694 16522
tri 41694 16514 41702 16522 sw
tri 41426 16506 41434 16514 ne
rect 41434 16506 41702 16514
tri 41702 16506 41710 16514 sw
rect 70802 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41434 16498 41442 16506 ne
rect 41442 16498 41710 16506
tri 41710 16498 41718 16506 sw
tri 41442 16490 41450 16498 ne
rect 41450 16490 41718 16498
tri 41718 16490 41726 16498 sw
tri 41450 16482 41458 16490 ne
rect 41458 16482 41726 16490
tri 41726 16482 41734 16490 sw
tri 41458 16474 41466 16482 ne
rect 41466 16474 41734 16482
tri 41734 16474 41742 16482 sw
tri 41466 16466 41474 16474 ne
rect 41474 16466 41742 16474
tri 41742 16466 41750 16474 sw
tri 41474 16458 41482 16466 ne
rect 41482 16458 41750 16466
tri 41750 16458 41758 16466 sw
tri 41482 16450 41490 16458 ne
rect 41490 16454 41758 16458
tri 41758 16454 41762 16458 sw
rect 41490 16450 41762 16454
tri 41762 16450 41766 16454 sw
rect 70802 16452 71000 16510
tri 41490 16442 41498 16450 ne
rect 41498 16444 41766 16450
rect 41498 16442 41634 16444
tri 41498 16438 41502 16442 ne
rect 41502 16438 41634 16442
tri 41502 16434 41506 16438 ne
rect 41506 16434 41634 16438
tri 41506 16426 41514 16434 ne
rect 41514 16426 41634 16434
tri 41514 16418 41522 16426 ne
rect 41522 16418 41634 16426
tri 41522 16410 41530 16418 ne
rect 41530 16410 41634 16418
tri 41530 16402 41538 16410 ne
rect 41538 16402 41634 16410
tri 41538 16394 41546 16402 ne
rect 41546 16398 41634 16402
rect 41680 16442 41766 16444
tri 41766 16442 41774 16450 sw
rect 41680 16434 41774 16442
tri 41774 16434 41782 16442 sw
rect 41680 16426 41782 16434
tri 41782 16426 41790 16434 sw
rect 41680 16418 41790 16426
tri 41790 16418 41798 16426 sw
rect 41680 16410 41798 16418
tri 41798 16410 41806 16418 sw
rect 41680 16402 41806 16410
tri 41806 16402 41814 16410 sw
rect 70802 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 41680 16398 41814 16402
rect 41546 16394 41814 16398
tri 41814 16394 41822 16402 sw
tri 41546 16386 41554 16394 ne
rect 41554 16386 41822 16394
tri 41822 16386 41830 16394 sw
tri 41554 16378 41562 16386 ne
rect 41562 16378 41830 16386
tri 41830 16378 41838 16386 sw
tri 41562 16370 41570 16378 ne
rect 41570 16370 41838 16378
tri 41838 16370 41846 16378 sw
tri 41570 16362 41578 16370 ne
rect 41578 16362 41846 16370
tri 41846 16362 41854 16370 sw
tri 41578 16354 41586 16362 ne
rect 41586 16354 41854 16362
tri 41854 16354 41862 16362 sw
tri 41586 16346 41594 16354 ne
rect 41594 16346 41862 16354
tri 41862 16346 41870 16354 sw
rect 70802 16348 71000 16406
tri 41594 16338 41602 16346 ne
rect 41602 16338 41870 16346
tri 41870 16338 41878 16346 sw
tri 41602 16330 41610 16338 ne
rect 41610 16330 41878 16338
tri 41878 16330 41886 16338 sw
tri 41610 16322 41618 16330 ne
rect 41618 16322 41886 16330
tri 41886 16322 41894 16330 sw
tri 41618 16314 41626 16322 ne
rect 41626 16314 41894 16322
tri 41894 16314 41902 16322 sw
tri 41626 16306 41634 16314 ne
rect 41634 16312 41902 16314
rect 41634 16306 41766 16312
tri 41634 16298 41642 16306 ne
rect 41642 16298 41766 16306
tri 41642 16290 41650 16298 ne
rect 41650 16290 41766 16298
tri 41650 16282 41658 16290 ne
rect 41658 16282 41766 16290
tri 41658 16274 41666 16282 ne
rect 41666 16274 41766 16282
tri 41666 16266 41674 16274 ne
rect 41674 16266 41766 16274
rect 41812 16306 41902 16312
tri 41902 16306 41910 16314 sw
rect 41812 16298 41910 16306
tri 41910 16298 41918 16306 sw
rect 70802 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16290 41918 16298
tri 41918 16290 41926 16298 sw
rect 41812 16282 41926 16290
tri 41926 16282 41934 16290 sw
rect 41812 16274 41934 16282
tri 41934 16274 41942 16282 sw
rect 41812 16266 41942 16274
tri 41942 16266 41950 16274 sw
tri 41674 16258 41682 16266 ne
rect 41682 16258 41950 16266
tri 41950 16258 41958 16266 sw
tri 41682 16250 41690 16258 ne
rect 41690 16250 41958 16258
tri 41958 16250 41966 16258 sw
tri 41690 16242 41698 16250 ne
rect 41698 16243 41966 16250
tri 41966 16243 41973 16250 sw
rect 70802 16244 71000 16302
rect 41698 16242 41973 16243
tri 41698 16234 41706 16242 ne
rect 41706 16235 41973 16242
tri 41973 16235 41981 16243 sw
rect 41706 16234 41981 16235
tri 41706 16226 41714 16234 ne
rect 41714 16227 41981 16234
tri 41981 16227 41989 16235 sw
rect 41714 16226 41989 16227
tri 41714 16218 41722 16226 ne
rect 41722 16219 41989 16226
tri 41989 16219 41997 16227 sw
rect 41722 16218 41997 16219
tri 41722 16210 41730 16218 ne
rect 41730 16211 41997 16218
tri 41997 16211 42005 16219 sw
rect 41730 16210 42005 16211
tri 41730 16202 41738 16210 ne
rect 41738 16203 42005 16210
tri 42005 16203 42013 16211 sw
rect 41738 16202 42013 16203
tri 41738 16194 41746 16202 ne
rect 41746 16195 42013 16202
tri 42013 16195 42021 16203 sw
rect 70802 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 41746 16194 42021 16195
tri 41746 16186 41754 16194 ne
rect 41754 16187 42021 16194
tri 42021 16187 42029 16195 sw
rect 41754 16186 42029 16187
tri 41754 16178 41762 16186 ne
rect 41762 16180 42029 16186
rect 41762 16178 41898 16180
tri 41762 16170 41770 16178 ne
rect 41770 16170 41898 16178
tri 41770 16162 41778 16170 ne
rect 41778 16162 41898 16170
tri 41778 16154 41786 16162 ne
rect 41786 16154 41898 16162
tri 41786 16146 41794 16154 ne
rect 41794 16146 41898 16154
tri 41794 16138 41802 16146 ne
rect 41802 16138 41898 16146
tri 41802 16130 41810 16138 ne
rect 41810 16134 41898 16138
rect 41944 16179 42029 16180
tri 42029 16179 42037 16187 sw
rect 41944 16171 42037 16179
tri 42037 16171 42045 16179 sw
rect 41944 16163 42045 16171
tri 42045 16163 42053 16171 sw
rect 41944 16155 42053 16163
tri 42053 16155 42061 16163 sw
rect 41944 16147 42061 16155
tri 42061 16147 42069 16155 sw
rect 41944 16139 42069 16147
tri 42069 16139 42077 16147 sw
rect 70802 16140 71000 16198
rect 41944 16134 42077 16139
rect 41810 16131 42077 16134
tri 42077 16131 42085 16139 sw
rect 41810 16130 42085 16131
tri 41810 16122 41818 16130 ne
rect 41818 16123 42085 16130
tri 42085 16123 42093 16131 sw
rect 41818 16122 42093 16123
tri 41818 16114 41826 16122 ne
rect 41826 16115 42093 16122
tri 42093 16115 42101 16123 sw
rect 41826 16114 42101 16115
tri 41826 16106 41834 16114 ne
rect 41834 16107 42101 16114
tri 42101 16107 42109 16115 sw
rect 41834 16106 42109 16107
tri 41834 16099 41841 16106 ne
rect 41841 16099 42109 16106
tri 42109 16099 42117 16107 sw
tri 41841 16091 41849 16099 ne
rect 41849 16091 42117 16099
tri 42117 16091 42125 16099 sw
rect 70802 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41849 16083 41857 16091 ne
rect 41857 16083 42125 16091
tri 42125 16083 42133 16091 sw
tri 41857 16075 41865 16083 ne
rect 41865 16075 42133 16083
tri 42133 16075 42141 16083 sw
tri 41865 16067 41873 16075 ne
rect 41873 16067 42141 16075
tri 42141 16067 42149 16075 sw
tri 41873 16059 41881 16067 ne
rect 41881 16059 42149 16067
tri 42149 16059 42157 16067 sw
tri 41881 16051 41889 16059 ne
rect 41889 16051 42157 16059
tri 42157 16051 42165 16059 sw
tri 41889 16043 41897 16051 ne
rect 41897 16048 42165 16051
rect 41897 16043 42030 16048
tri 41897 16035 41905 16043 ne
rect 41905 16035 42030 16043
tri 41905 16027 41913 16035 ne
rect 41913 16027 42030 16035
tri 41913 16019 41921 16027 ne
rect 41921 16019 42030 16027
tri 41921 16011 41929 16019 ne
rect 41929 16011 42030 16019
tri 41929 16003 41937 16011 ne
rect 41937 16003 42030 16011
tri 41937 15995 41945 16003 ne
rect 41945 16002 42030 16003
rect 42076 16043 42165 16048
tri 42165 16043 42173 16051 sw
rect 42076 16035 42173 16043
tri 42173 16035 42181 16043 sw
rect 70802 16036 71000 16094
rect 42076 16027 42181 16035
tri 42181 16027 42189 16035 sw
rect 42076 16019 42189 16027
tri 42189 16019 42197 16027 sw
rect 42076 16015 42197 16019
tri 42197 16015 42201 16019 sw
rect 42076 16007 42201 16015
tri 42201 16007 42209 16015 sw
rect 42076 16002 42209 16007
rect 41945 15999 42209 16002
tri 42209 15999 42217 16007 sw
rect 41945 15995 42217 15999
tri 41945 15987 41953 15995 ne
rect 41953 15991 42217 15995
tri 42217 15991 42225 15999 sw
rect 41953 15987 42225 15991
tri 41953 15979 41961 15987 ne
rect 41961 15983 42225 15987
tri 42225 15983 42233 15991 sw
rect 70802 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
rect 41961 15979 42233 15983
tri 41961 15978 41962 15979 ne
rect 41962 15978 42233 15979
tri 41962 15970 41970 15978 ne
rect 41970 15975 42233 15978
tri 42233 15975 42241 15983 sw
rect 41970 15970 42241 15975
tri 41970 15962 41978 15970 ne
rect 41978 15967 42241 15970
tri 42241 15967 42249 15975 sw
rect 41978 15962 42249 15967
tri 41978 15954 41986 15962 ne
rect 41986 15959 42249 15962
tri 42249 15959 42257 15967 sw
rect 41986 15954 42257 15959
tri 41986 15946 41994 15954 ne
rect 41994 15951 42257 15954
tri 42257 15951 42265 15959 sw
rect 41994 15946 42265 15951
tri 41994 15938 42002 15946 ne
rect 42002 15943 42265 15946
tri 42265 15943 42273 15951 sw
rect 42002 15938 42273 15943
tri 42002 15930 42010 15938 ne
rect 42010 15935 42273 15938
tri 42273 15935 42281 15943 sw
rect 42010 15930 42281 15935
tri 42010 15922 42018 15930 ne
rect 42018 15927 42281 15930
tri 42281 15927 42289 15935 sw
rect 70802 15932 71000 15990
rect 42018 15922 42289 15927
tri 42289 15922 42294 15927 sw
tri 42018 15914 42026 15922 ne
rect 42026 15916 42294 15922
rect 42026 15914 42162 15916
tri 42026 15906 42034 15914 ne
rect 42034 15906 42162 15914
tri 42034 15898 42042 15906 ne
rect 42042 15898 42162 15906
tri 42042 15890 42050 15898 ne
rect 42050 15890 42162 15898
tri 42050 15882 42058 15890 ne
rect 42058 15882 42162 15890
tri 42058 15874 42066 15882 ne
rect 42066 15874 42162 15882
tri 42066 15866 42074 15874 ne
rect 42074 15870 42162 15874
rect 42208 15914 42294 15916
tri 42294 15914 42302 15922 sw
rect 42208 15906 42302 15914
tri 42302 15906 42310 15914 sw
rect 42208 15898 42310 15906
tri 42310 15898 42318 15906 sw
rect 42208 15890 42318 15898
tri 42318 15890 42326 15898 sw
rect 42208 15882 42326 15890
tri 42326 15882 42334 15890 sw
rect 70802 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 42208 15874 42334 15882
tri 42334 15874 42342 15882 sw
rect 42208 15870 42342 15874
rect 42074 15866 42342 15870
tri 42342 15866 42350 15874 sw
tri 42074 15858 42082 15866 ne
rect 42082 15860 42350 15866
tri 42350 15860 42356 15866 sw
rect 42082 15858 42356 15860
tri 42082 15852 42088 15858 ne
rect 42088 15852 42356 15858
tri 42356 15852 42364 15860 sw
tri 42088 15844 42096 15852 ne
rect 42096 15844 42364 15852
tri 42364 15844 42372 15852 sw
tri 42096 15836 42104 15844 ne
rect 42104 15836 42372 15844
tri 42372 15836 42380 15844 sw
tri 42104 15828 42112 15836 ne
rect 42112 15828 42380 15836
tri 42380 15828 42388 15836 sw
rect 70802 15828 71000 15886
tri 42112 15820 42120 15828 ne
rect 42120 15820 42388 15828
tri 42388 15820 42396 15828 sw
tri 42120 15812 42128 15820 ne
rect 42128 15812 42396 15820
tri 42396 15812 42404 15820 sw
tri 42128 15804 42136 15812 ne
rect 42136 15804 42404 15812
tri 42404 15804 42412 15812 sw
tri 42136 15796 42144 15804 ne
rect 42144 15796 42412 15804
tri 42412 15796 42420 15804 sw
tri 42144 15788 42152 15796 ne
rect 42152 15788 42420 15796
tri 42420 15788 42428 15796 sw
tri 42152 15780 42160 15788 ne
rect 42160 15784 42428 15788
rect 42160 15780 42294 15784
tri 42160 15772 42168 15780 ne
rect 42168 15772 42294 15780
tri 42168 15764 42176 15772 ne
rect 42176 15764 42294 15772
tri 42176 15756 42184 15764 ne
rect 42184 15756 42294 15764
tri 42184 15748 42192 15756 ne
rect 42192 15748 42294 15756
tri 42192 15740 42200 15748 ne
rect 42200 15740 42294 15748
tri 42200 15739 42201 15740 ne
rect 42201 15739 42294 15740
tri 42201 15731 42209 15739 ne
rect 42209 15738 42294 15739
rect 42340 15780 42428 15784
tri 42428 15780 42436 15788 sw
rect 70802 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15772 42436 15780
tri 42436 15772 42444 15780 sw
rect 42340 15764 42444 15772
tri 42444 15764 42452 15772 sw
rect 42340 15756 42452 15764
tri 42452 15756 42460 15764 sw
rect 42340 15748 42460 15756
tri 42460 15748 42468 15756 sw
rect 42340 15744 42468 15748
tri 42468 15744 42472 15748 sw
rect 42340 15738 42472 15744
rect 42209 15736 42472 15738
tri 42472 15736 42480 15744 sw
rect 42209 15731 42480 15736
tri 42209 15723 42217 15731 ne
rect 42217 15728 42480 15731
tri 42480 15728 42488 15736 sw
rect 42217 15723 42488 15728
tri 42217 15715 42225 15723 ne
rect 42225 15720 42488 15723
tri 42488 15720 42496 15728 sw
rect 70802 15724 71000 15782
rect 42225 15715 42496 15720
tri 42225 15707 42233 15715 ne
rect 42233 15712 42496 15715
tri 42496 15712 42504 15720 sw
rect 42233 15707 42504 15712
tri 42233 15699 42241 15707 ne
rect 42241 15704 42504 15707
tri 42504 15704 42512 15712 sw
rect 42241 15699 42512 15704
tri 42241 15691 42249 15699 ne
rect 42249 15696 42512 15699
tri 42512 15696 42520 15704 sw
rect 42249 15691 42520 15696
tri 42249 15683 42257 15691 ne
rect 42257 15688 42520 15691
tri 42520 15688 42528 15696 sw
rect 42257 15683 42528 15688
tri 42257 15675 42265 15683 ne
rect 42265 15680 42528 15683
tri 42528 15680 42536 15688 sw
rect 42265 15675 42536 15680
tri 42265 15667 42273 15675 ne
rect 42273 15672 42536 15675
tri 42536 15672 42544 15680 sw
rect 70802 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
rect 42273 15667 42544 15672
tri 42544 15667 42549 15672 sw
tri 42273 15659 42281 15667 ne
rect 42281 15659 42549 15667
tri 42549 15659 42557 15667 sw
tri 42281 15651 42289 15659 ne
rect 42289 15652 42557 15659
rect 42289 15651 42426 15652
tri 42289 15643 42297 15651 ne
rect 42297 15643 42426 15651
tri 42297 15635 42305 15643 ne
rect 42305 15635 42426 15643
tri 42305 15627 42313 15635 ne
rect 42313 15627 42426 15635
tri 42313 15619 42321 15627 ne
rect 42321 15619 42426 15627
tri 42321 15611 42329 15619 ne
rect 42329 15611 42426 15619
tri 42329 15605 42335 15611 ne
rect 42335 15606 42426 15611
rect 42472 15651 42557 15652
tri 42557 15651 42565 15659 sw
rect 42472 15643 42565 15651
tri 42565 15643 42573 15651 sw
rect 42472 15635 42573 15643
tri 42573 15635 42581 15643 sw
rect 42472 15627 42581 15635
tri 42581 15627 42589 15635 sw
rect 42472 15619 42589 15627
tri 42589 15619 42597 15627 sw
rect 70802 15620 71000 15678
rect 42472 15611 42597 15619
tri 42597 15611 42605 15619 sw
rect 42472 15606 42605 15611
rect 42335 15605 42605 15606
tri 42335 15597 42343 15605 ne
rect 42343 15603 42605 15605
tri 42605 15603 42613 15611 sw
rect 42343 15597 42613 15603
tri 42343 15589 42351 15597 ne
rect 42351 15595 42613 15597
tri 42613 15595 42621 15603 sw
rect 42351 15592 42621 15595
tri 42621 15592 42624 15595 sw
rect 42351 15589 42624 15592
tri 42351 15581 42359 15589 ne
rect 42359 15584 42624 15589
tri 42624 15584 42632 15592 sw
rect 42359 15581 42632 15584
tri 42359 15573 42367 15581 ne
rect 42367 15576 42632 15581
tri 42632 15576 42640 15584 sw
rect 42367 15573 42640 15576
tri 42367 15565 42375 15573 ne
rect 42375 15568 42640 15573
tri 42640 15568 42648 15576 sw
rect 70802 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
rect 42375 15565 42648 15568
tri 42375 15557 42383 15565 ne
rect 42383 15560 42648 15565
tri 42648 15560 42656 15568 sw
rect 42383 15557 42656 15560
tri 42383 15549 42391 15557 ne
rect 42391 15552 42656 15557
tri 42656 15552 42664 15560 sw
rect 42391 15549 42664 15552
tri 42391 15541 42399 15549 ne
rect 42399 15544 42664 15549
tri 42664 15544 42672 15552 sw
rect 42399 15541 42672 15544
tri 42399 15533 42407 15541 ne
rect 42407 15536 42672 15541
tri 42672 15536 42680 15544 sw
rect 42407 15533 42680 15536
tri 42407 15525 42415 15533 ne
rect 42415 15528 42680 15533
tri 42680 15528 42688 15536 sw
rect 42415 15525 42688 15528
tri 42415 15517 42423 15525 ne
rect 42423 15520 42688 15525
tri 42688 15520 42696 15528 sw
rect 42423 15517 42558 15520
tri 42423 15509 42431 15517 ne
rect 42431 15509 42558 15517
tri 42431 15501 42439 15509 ne
rect 42439 15501 42558 15509
tri 42439 15493 42447 15501 ne
rect 42447 15493 42558 15501
tri 42447 15485 42455 15493 ne
rect 42455 15485 42558 15493
tri 42455 15477 42463 15485 ne
rect 42463 15477 42558 15485
tri 42463 15472 42468 15477 ne
rect 42468 15474 42558 15477
rect 42604 15512 42696 15520
tri 42696 15512 42704 15520 sw
rect 70802 15516 71000 15574
rect 42604 15504 42704 15512
tri 42704 15504 42712 15512 sw
rect 42604 15496 42712 15504
tri 42712 15496 42720 15504 sw
rect 42604 15488 42720 15496
tri 42720 15488 42728 15496 sw
rect 42604 15480 42728 15488
tri 42728 15480 42736 15488 sw
rect 42604 15474 42736 15480
rect 42468 15472 42736 15474
tri 42736 15472 42744 15480 sw
tri 42468 15464 42476 15472 ne
rect 42476 15471 42744 15472
tri 42744 15471 42745 15472 sw
rect 42476 15464 42745 15471
tri 42476 15456 42484 15464 ne
rect 42484 15463 42745 15464
tri 42745 15463 42753 15471 sw
rect 70802 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 42484 15456 42753 15463
tri 42484 15448 42492 15456 ne
rect 42492 15455 42753 15456
tri 42753 15455 42761 15463 sw
rect 42492 15448 42761 15455
tri 42492 15440 42500 15448 ne
rect 42500 15447 42761 15448
tri 42761 15447 42769 15455 sw
rect 42500 15440 42769 15447
tri 42500 15432 42508 15440 ne
rect 42508 15439 42769 15440
tri 42769 15439 42777 15447 sw
rect 42508 15432 42777 15439
tri 42508 15424 42516 15432 ne
rect 42516 15431 42777 15432
tri 42777 15431 42785 15439 sw
rect 42516 15424 42785 15431
tri 42516 15416 42524 15424 ne
rect 42524 15423 42785 15424
tri 42785 15423 42793 15431 sw
rect 42524 15416 42793 15423
tri 42524 15408 42532 15416 ne
rect 42532 15415 42793 15416
tri 42793 15415 42801 15423 sw
rect 42532 15408 42801 15415
tri 42532 15400 42540 15408 ne
rect 42540 15407 42801 15408
tri 42801 15407 42809 15415 sw
rect 70802 15412 71000 15470
rect 42540 15400 42809 15407
tri 42540 15396 42544 15400 ne
rect 42544 15399 42809 15400
tri 42809 15399 42817 15407 sw
rect 42544 15396 42817 15399
tri 42544 15392 42548 15396 ne
rect 42548 15392 42817 15396
tri 42817 15392 42824 15399 sw
tri 42548 15384 42556 15392 ne
rect 42556 15391 42824 15392
tri 42824 15391 42825 15392 sw
rect 42556 15388 42825 15391
rect 42556 15384 42690 15388
tri 42556 15376 42564 15384 ne
rect 42564 15376 42690 15384
tri 42564 15368 42572 15376 ne
rect 42572 15368 42690 15376
tri 42572 15360 42580 15368 ne
rect 42580 15360 42690 15368
tri 42580 15352 42588 15360 ne
rect 42588 15352 42690 15360
tri 42588 15344 42596 15352 ne
rect 42596 15344 42690 15352
tri 42596 15336 42604 15344 ne
rect 42604 15342 42690 15344
rect 42736 15383 42825 15388
tri 42825 15383 42833 15391 sw
rect 42736 15375 42833 15383
tri 42833 15375 42841 15383 sw
rect 42736 15367 42841 15375
tri 42841 15367 42849 15375 sw
rect 42736 15359 42849 15367
tri 42849 15359 42857 15367 sw
rect 70802 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15351 42857 15359
tri 42857 15351 42865 15359 sw
rect 42736 15343 42865 15351
tri 42865 15343 42873 15351 sw
rect 42736 15342 42873 15343
rect 42604 15336 42873 15342
tri 42604 15328 42612 15336 ne
rect 42612 15335 42873 15336
tri 42873 15335 42881 15343 sw
rect 42612 15328 42881 15335
tri 42612 15325 42615 15328 ne
rect 42615 15327 42881 15328
tri 42881 15327 42889 15335 sw
rect 42615 15325 42889 15327
tri 42889 15325 42891 15327 sw
tri 42615 15317 42623 15325 ne
rect 42623 15317 42891 15325
tri 42891 15317 42899 15325 sw
tri 42623 15309 42631 15317 ne
rect 42631 15309 42899 15317
tri 42899 15309 42907 15317 sw
tri 42631 15301 42639 15309 ne
rect 42639 15301 42907 15309
tri 42907 15301 42915 15309 sw
rect 70802 15308 71000 15366
tri 42639 15293 42647 15301 ne
rect 42647 15293 42915 15301
tri 42915 15293 42923 15301 sw
tri 42647 15285 42655 15293 ne
rect 42655 15285 42923 15293
tri 42923 15285 42931 15293 sw
tri 42655 15277 42663 15285 ne
rect 42663 15277 42931 15285
tri 42931 15277 42939 15285 sw
tri 42663 15269 42671 15277 ne
rect 42671 15269 42939 15277
tri 42939 15269 42947 15277 sw
tri 42671 15261 42679 15269 ne
rect 42679 15261 42947 15269
tri 42947 15261 42955 15269 sw
rect 70802 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
tri 42679 15253 42687 15261 ne
rect 42687 15256 42955 15261
rect 42687 15253 42822 15256
tri 42687 15245 42695 15253 ne
rect 42695 15245 42822 15253
tri 42695 15237 42703 15245 ne
rect 42703 15237 42822 15245
tri 42703 15229 42711 15237 ne
rect 42711 15229 42822 15237
tri 42711 15221 42719 15229 ne
rect 42719 15221 42822 15229
tri 42719 15213 42727 15221 ne
rect 42727 15213 42822 15221
tri 42727 15205 42735 15213 ne
rect 42735 15210 42822 15213
rect 42868 15253 42955 15256
tri 42955 15253 42963 15261 sw
rect 42868 15245 42963 15253
tri 42963 15245 42971 15253 sw
rect 42868 15237 42971 15245
tri 42971 15237 42979 15245 sw
rect 42868 15229 42979 15237
tri 42979 15229 42987 15237 sw
rect 42868 15221 42987 15229
tri 42987 15221 42995 15229 sw
rect 42868 15213 42995 15221
tri 42995 15213 43003 15221 sw
rect 42868 15210 43003 15213
rect 42735 15205 43003 15210
tri 43003 15205 43011 15213 sw
tri 42735 15197 42743 15205 ne
rect 42743 15197 43011 15205
tri 43011 15197 43019 15205 sw
rect 70802 15204 71000 15262
tri 42743 15189 42751 15197 ne
rect 42751 15191 43019 15197
tri 43019 15191 43025 15197 sw
rect 42751 15189 43025 15191
tri 42751 15186 42754 15189 ne
rect 42754 15186 43025 15189
tri 42754 15178 42762 15186 ne
rect 42762 15183 43025 15186
tri 43025 15183 43033 15191 sw
rect 42762 15178 43033 15183
tri 42762 15170 42770 15178 ne
rect 42770 15175 43033 15178
tri 43033 15175 43041 15183 sw
rect 42770 15170 43041 15175
tri 42770 15162 42778 15170 ne
rect 42778 15167 43041 15170
tri 43041 15167 43049 15175 sw
rect 42778 15162 43049 15167
tri 42778 15154 42786 15162 ne
rect 42786 15159 43049 15162
tri 43049 15159 43057 15167 sw
rect 42786 15154 43057 15159
tri 42786 15146 42794 15154 ne
rect 42794 15151 43057 15154
tri 43057 15151 43065 15159 sw
rect 70802 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
rect 42794 15146 43065 15151
tri 42794 15138 42802 15146 ne
rect 42802 15143 43065 15146
tri 43065 15143 43073 15151 sw
rect 42802 15138 43073 15143
tri 42802 15130 42810 15138 ne
rect 42810 15135 43073 15138
tri 43073 15135 43081 15143 sw
rect 42810 15130 43081 15135
tri 42810 15122 42818 15130 ne
rect 42818 15127 43081 15130
tri 43081 15127 43089 15135 sw
rect 42818 15124 43089 15127
rect 42818 15122 42954 15124
tri 42818 15119 42821 15122 ne
rect 42821 15119 42954 15122
tri 42821 15114 42826 15119 ne
rect 42826 15114 42954 15119
tri 42826 15106 42834 15114 ne
rect 42834 15106 42954 15114
tri 42834 15098 42842 15106 ne
rect 42842 15098 42954 15106
tri 42842 15090 42850 15098 ne
rect 42850 15090 42954 15098
tri 42850 15082 42858 15090 ne
rect 42858 15082 42954 15090
tri 42858 15074 42866 15082 ne
rect 42866 15078 42954 15082
rect 43000 15119 43089 15124
tri 43089 15119 43097 15127 sw
rect 43000 15114 43097 15119
tri 43097 15114 43102 15119 sw
rect 43000 15111 43102 15114
tri 43102 15111 43105 15114 sw
rect 43000 15103 43105 15111
tri 43105 15103 43113 15111 sw
rect 43000 15095 43113 15103
tri 43113 15095 43121 15103 sw
rect 70802 15100 71000 15158
rect 43000 15087 43121 15095
tri 43121 15087 43129 15095 sw
rect 43000 15079 43129 15087
tri 43129 15079 43137 15087 sw
rect 43000 15078 43137 15079
rect 42866 15074 43137 15078
tri 42866 15069 42871 15074 ne
rect 42871 15071 43137 15074
tri 43137 15071 43145 15079 sw
rect 42871 15069 43145 15071
tri 43145 15069 43147 15071 sw
tri 42871 15061 42879 15069 ne
rect 42879 15061 43147 15069
tri 43147 15061 43155 15069 sw
tri 42879 15053 42887 15061 ne
rect 42887 15053 43155 15061
tri 43155 15053 43163 15061 sw
rect 70802 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42887 15045 42895 15053 ne
rect 42895 15045 43163 15053
tri 43163 15045 43171 15053 sw
tri 42895 15037 42903 15045 ne
rect 42903 15037 43171 15045
tri 43171 15037 43179 15045 sw
tri 42903 15029 42911 15037 ne
rect 42911 15029 43179 15037
tri 43179 15029 43187 15037 sw
tri 42911 15021 42919 15029 ne
rect 42919 15021 43187 15029
tri 43187 15021 43195 15029 sw
tri 42919 15013 42927 15021 ne
rect 42927 15013 43195 15021
tri 43195 15013 43203 15021 sw
tri 42927 15005 42935 15013 ne
rect 42935 15005 43203 15013
tri 43203 15005 43211 15013 sw
tri 42935 14997 42943 15005 ne
rect 42943 14997 43211 15005
tri 43211 14997 43219 15005 sw
tri 42943 14989 42951 14997 ne
rect 42951 14992 43219 14997
rect 42951 14989 43086 14992
tri 42951 14981 42959 14989 ne
rect 42959 14981 43086 14989
tri 42959 14973 42967 14981 ne
rect 42967 14973 43086 14981
tri 42967 14965 42975 14973 ne
rect 42975 14965 43086 14973
tri 42975 14957 42983 14965 ne
rect 42983 14957 43086 14965
tri 42983 14949 42991 14957 ne
rect 42991 14949 43086 14957
tri 42991 14941 42999 14949 ne
rect 42999 14946 43086 14949
rect 43132 14989 43219 14992
tri 43219 14989 43227 14997 sw
rect 70802 14996 71000 15054
rect 43132 14981 43227 14989
tri 43227 14981 43235 14989 sw
rect 43132 14973 43235 14981
tri 43235 14973 43243 14981 sw
rect 43132 14965 43243 14973
tri 43243 14965 43251 14973 sw
rect 43132 14957 43251 14965
tri 43251 14957 43259 14965 sw
rect 43132 14949 43259 14957
tri 43259 14949 43267 14957 sw
rect 70802 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 43132 14946 43267 14949
rect 42999 14941 43267 14946
tri 43267 14941 43275 14949 sw
tri 42999 14933 43007 14941 ne
rect 43007 14933 43275 14941
tri 43275 14933 43283 14941 sw
tri 43007 14931 43009 14933 ne
rect 43009 14931 43283 14933
tri 43283 14931 43285 14933 sw
tri 43009 14923 43017 14931 ne
rect 43017 14923 43285 14931
tri 43285 14923 43293 14931 sw
tri 43017 14915 43025 14923 ne
rect 43025 14915 43293 14923
tri 43293 14915 43301 14923 sw
tri 43025 14907 43033 14915 ne
rect 43033 14907 43301 14915
tri 43301 14907 43309 14915 sw
tri 43033 14899 43041 14907 ne
rect 43041 14899 43309 14907
tri 43309 14899 43317 14907 sw
tri 43041 14891 43049 14899 ne
rect 43049 14891 43317 14899
tri 43317 14891 43325 14899 sw
rect 70802 14892 71000 14950
tri 43049 14883 43057 14891 ne
rect 43057 14883 43325 14891
tri 43325 14883 43333 14891 sw
tri 43057 14875 43065 14883 ne
rect 43065 14875 43333 14883
tri 43333 14875 43341 14883 sw
tri 43065 14867 43073 14875 ne
rect 43073 14867 43341 14875
tri 43341 14867 43349 14875 sw
tri 43073 14859 43081 14867 ne
rect 43081 14860 43349 14867
rect 43081 14859 43218 14860
tri 43081 14851 43089 14859 ne
rect 43089 14851 43218 14859
tri 43089 14843 43097 14851 ne
rect 43097 14843 43218 14851
tri 43097 14835 43105 14843 ne
rect 43105 14835 43218 14843
tri 43105 14827 43113 14835 ne
rect 43113 14827 43218 14835
tri 43113 14819 43121 14827 ne
rect 43121 14819 43218 14827
tri 43121 14811 43129 14819 ne
rect 43129 14814 43218 14819
rect 43264 14859 43349 14860
tri 43349 14859 43357 14867 sw
rect 43264 14851 43357 14859
tri 43357 14851 43365 14859 sw
rect 43264 14843 43365 14851
tri 43365 14843 43373 14851 sw
rect 70802 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 43264 14835 43373 14843
tri 43373 14835 43381 14843 sw
rect 43264 14827 43381 14835
tri 43381 14827 43389 14835 sw
rect 43264 14819 43389 14827
tri 43389 14819 43397 14827 sw
rect 43264 14814 43397 14819
rect 43129 14811 43397 14814
tri 43397 14811 43405 14819 sw
tri 43129 14803 43137 14811 ne
rect 43137 14803 43405 14811
tri 43405 14803 43413 14811 sw
tri 43137 14795 43145 14803 ne
rect 43145 14795 43413 14803
tri 43413 14795 43421 14803 sw
tri 43145 14787 43153 14795 ne
rect 43153 14787 43421 14795
tri 43421 14787 43429 14795 sw
rect 70802 14788 71000 14846
tri 43153 14785 43155 14787 ne
rect 43155 14785 43429 14787
tri 43429 14785 43431 14787 sw
tri 43155 14777 43163 14785 ne
rect 43163 14777 43431 14785
tri 43431 14777 43439 14785 sw
tri 43163 14769 43171 14777 ne
rect 43171 14769 43439 14777
tri 43439 14769 43447 14777 sw
tri 43171 14761 43179 14769 ne
rect 43179 14761 43447 14769
tri 43447 14761 43455 14769 sw
tri 43179 14753 43187 14761 ne
rect 43187 14753 43455 14761
tri 43455 14753 43463 14761 sw
tri 43187 14745 43195 14753 ne
rect 43195 14745 43463 14753
tri 43463 14745 43471 14753 sw
tri 43195 14737 43203 14745 ne
rect 43203 14737 43471 14745
tri 43471 14737 43479 14745 sw
rect 70802 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
tri 43203 14729 43211 14737 ne
rect 43211 14729 43479 14737
tri 43479 14729 43487 14737 sw
tri 43211 14721 43219 14729 ne
rect 43219 14728 43487 14729
rect 43219 14721 43350 14728
tri 43219 14713 43227 14721 ne
rect 43227 14713 43350 14721
tri 43227 14705 43235 14713 ne
rect 43235 14705 43350 14713
tri 43235 14697 43243 14705 ne
rect 43243 14697 43350 14705
tri 43243 14689 43251 14697 ne
rect 43251 14689 43350 14697
tri 43251 14681 43259 14689 ne
rect 43259 14682 43350 14689
rect 43396 14721 43487 14728
tri 43487 14721 43495 14729 sw
rect 43396 14713 43495 14721
tri 43495 14713 43503 14721 sw
rect 43396 14705 43503 14713
tri 43503 14705 43511 14713 sw
rect 43396 14697 43511 14705
tri 43511 14697 43519 14705 sw
rect 43396 14689 43519 14697
tri 43519 14689 43527 14697 sw
rect 43396 14683 43527 14689
tri 43527 14683 43533 14689 sw
rect 70802 14684 71000 14742
rect 43396 14682 43533 14683
rect 43259 14681 43533 14682
tri 43259 14673 43267 14681 ne
rect 43267 14675 43533 14681
tri 43533 14675 43541 14683 sw
rect 43267 14673 43541 14675
tri 43267 14666 43274 14673 ne
rect 43274 14667 43541 14673
tri 43541 14667 43549 14675 sw
rect 43274 14666 43549 14667
tri 43274 14658 43282 14666 ne
rect 43282 14659 43549 14666
tri 43549 14659 43557 14667 sw
rect 43282 14658 43557 14659
tri 43282 14650 43290 14658 ne
rect 43290 14651 43557 14658
tri 43557 14651 43565 14659 sw
rect 43290 14650 43565 14651
tri 43290 14642 43298 14650 ne
rect 43298 14643 43565 14650
tri 43565 14643 43573 14651 sw
rect 43298 14642 43573 14643
tri 43298 14634 43306 14642 ne
rect 43306 14635 43573 14642
tri 43573 14635 43581 14643 sw
rect 70802 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
rect 43306 14634 43581 14635
tri 43306 14626 43314 14634 ne
rect 43314 14627 43581 14634
tri 43581 14627 43589 14635 sw
rect 43314 14626 43589 14627
tri 43314 14618 43322 14626 ne
rect 43322 14619 43589 14626
tri 43589 14619 43597 14627 sw
rect 43322 14618 43597 14619
tri 43322 14610 43330 14618 ne
rect 43330 14611 43597 14618
tri 43597 14611 43605 14619 sw
rect 43330 14610 43605 14611
tri 43330 14602 43338 14610 ne
rect 43338 14607 43605 14610
tri 43605 14607 43609 14611 sw
rect 43338 14602 43609 14607
tri 43338 14594 43346 14602 ne
rect 43346 14599 43609 14602
tri 43609 14599 43617 14607 sw
rect 43346 14596 43617 14599
rect 43346 14594 43482 14596
tri 43346 14590 43350 14594 ne
rect 43350 14590 43482 14594
tri 43350 14586 43354 14590 ne
rect 43354 14586 43482 14590
tri 43354 14578 43362 14586 ne
rect 43362 14578 43482 14586
tri 43362 14570 43370 14578 ne
rect 43370 14570 43482 14578
tri 43370 14562 43378 14570 ne
rect 43378 14562 43482 14570
tri 43378 14554 43386 14562 ne
rect 43386 14554 43482 14562
tri 43386 14546 43394 14554 ne
rect 43394 14550 43482 14554
rect 43528 14591 43617 14596
tri 43617 14591 43625 14599 sw
rect 43528 14586 43625 14591
tri 43625 14586 43630 14591 sw
rect 43528 14578 43630 14586
tri 43630 14578 43638 14586 sw
rect 70802 14580 71000 14638
rect 43528 14570 43638 14578
tri 43638 14570 43646 14578 sw
rect 43528 14562 43646 14570
tri 43646 14562 43654 14570 sw
rect 43528 14554 43654 14562
tri 43654 14554 43662 14562 sw
rect 43528 14550 43662 14554
rect 43394 14546 43662 14550
tri 43662 14546 43670 14554 sw
tri 43394 14538 43402 14546 ne
rect 43402 14538 43670 14546
tri 43670 14538 43678 14546 sw
tri 43402 14530 43410 14538 ne
rect 43410 14533 43678 14538
tri 43678 14533 43683 14538 sw
rect 70802 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
rect 43410 14530 43683 14533
tri 43410 14522 43418 14530 ne
rect 43418 14525 43683 14530
tri 43683 14525 43691 14533 sw
rect 43418 14522 43691 14525
tri 43418 14518 43422 14522 ne
rect 43422 14518 43691 14522
tri 43422 14510 43430 14518 ne
rect 43430 14517 43691 14518
tri 43691 14517 43699 14525 sw
rect 43430 14510 43699 14517
tri 43430 14502 43438 14510 ne
rect 43438 14509 43699 14510
tri 43699 14509 43707 14517 sw
rect 43438 14502 43707 14509
tri 43438 14494 43446 14502 ne
rect 43446 14501 43707 14502
tri 43707 14501 43715 14509 sw
rect 43446 14494 43715 14501
tri 43446 14486 43454 14494 ne
rect 43454 14493 43715 14494
tri 43715 14493 43723 14501 sw
rect 43454 14486 43723 14493
tri 43454 14478 43462 14486 ne
rect 43462 14485 43723 14486
tri 43723 14485 43731 14493 sw
rect 43462 14478 43731 14485
tri 43462 14470 43470 14478 ne
rect 43470 14477 43731 14478
tri 43731 14477 43739 14485 sw
rect 43470 14470 43739 14477
tri 43470 14462 43478 14470 ne
rect 43478 14469 43739 14470
tri 43739 14469 43747 14477 sw
rect 70802 14476 71000 14534
rect 43478 14464 43747 14469
rect 43478 14462 43614 14464
tri 43478 14454 43486 14462 ne
rect 43486 14454 43614 14462
tri 43486 14446 43494 14454 ne
rect 43494 14446 43614 14454
tri 43494 14438 43502 14446 ne
rect 43502 14438 43614 14446
tri 43502 14430 43510 14438 ne
rect 43510 14430 43614 14438
tri 43510 14422 43518 14430 ne
rect 43518 14422 43614 14430
tri 43518 14414 43526 14422 ne
rect 43526 14418 43614 14422
rect 43660 14461 43747 14464
tri 43747 14461 43755 14469 sw
rect 43660 14453 43755 14461
tri 43755 14453 43763 14461 sw
rect 43660 14445 43763 14453
tri 43763 14445 43771 14453 sw
rect 43660 14437 43771 14445
tri 43771 14437 43779 14445 sw
rect 43660 14429 43779 14437
tri 43779 14429 43787 14437 sw
rect 70802 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 43660 14421 43787 14429
tri 43787 14421 43795 14429 sw
rect 43660 14418 43795 14421
rect 43526 14414 43795 14418
tri 43526 14406 43534 14414 ne
rect 43534 14413 43795 14414
tri 43795 14413 43803 14421 sw
rect 43534 14406 43803 14413
tri 43534 14398 43542 14406 ne
rect 43542 14405 43803 14406
tri 43803 14405 43811 14413 sw
rect 43542 14398 43811 14405
tri 43542 14390 43550 14398 ne
rect 43550 14397 43811 14398
tri 43811 14397 43819 14405 sw
rect 43550 14395 43819 14397
tri 43819 14395 43821 14397 sw
rect 43550 14390 43821 14395
tri 43550 14387 43553 14390 ne
rect 43553 14387 43821 14390
tri 43821 14387 43829 14395 sw
tri 43553 14379 43561 14387 ne
rect 43561 14379 43829 14387
tri 43829 14379 43837 14387 sw
tri 43561 14371 43569 14379 ne
rect 43569 14371 43837 14379
tri 43837 14371 43845 14379 sw
rect 70802 14372 71000 14430
tri 43569 14363 43577 14371 ne
rect 43577 14363 43845 14371
tri 43845 14363 43853 14371 sw
tri 43577 14355 43585 14363 ne
rect 43585 14355 43853 14363
tri 43853 14355 43861 14363 sw
tri 43585 14347 43593 14355 ne
rect 43593 14347 43861 14355
tri 43861 14347 43869 14355 sw
tri 43593 14339 43601 14347 ne
rect 43601 14339 43869 14347
tri 43869 14339 43877 14347 sw
tri 43601 14331 43609 14339 ne
rect 43609 14332 43877 14339
rect 43609 14331 43746 14332
tri 43609 14323 43617 14331 ne
rect 43617 14323 43746 14331
tri 43617 14315 43625 14323 ne
rect 43625 14315 43746 14323
tri 43625 14307 43633 14315 ne
rect 43633 14307 43746 14315
tri 43633 14299 43641 14307 ne
rect 43641 14299 43746 14307
tri 43641 14291 43649 14299 ne
rect 43649 14291 43746 14299
tri 43649 14283 43657 14291 ne
rect 43657 14286 43746 14291
rect 43792 14331 43877 14332
tri 43877 14331 43885 14339 sw
rect 43792 14323 43885 14331
tri 43885 14323 43893 14331 sw
rect 70802 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43792 14315 43893 14323
tri 43893 14315 43901 14323 sw
rect 43792 14307 43901 14315
tri 43901 14307 43909 14315 sw
rect 43792 14299 43909 14307
tri 43909 14299 43917 14307 sw
rect 43792 14291 43917 14299
tri 43917 14291 43925 14299 sw
rect 43792 14286 43925 14291
rect 43657 14283 43925 14286
tri 43925 14283 43933 14291 sw
tri 43657 14275 43665 14283 ne
rect 43665 14275 43933 14283
tri 43933 14275 43941 14283 sw
tri 43665 14267 43673 14275 ne
rect 43673 14267 43941 14275
tri 43941 14267 43949 14275 sw
rect 70802 14268 71000 14326
tri 43673 14259 43681 14267 ne
rect 43681 14259 43949 14267
tri 43949 14259 43957 14267 sw
tri 43681 14251 43689 14259 ne
rect 43689 14251 43957 14259
tri 43957 14251 43965 14259 sw
tri 43689 14249 43691 14251 ne
rect 43691 14249 43965 14251
tri 43965 14249 43967 14251 sw
tri 43691 14241 43699 14249 ne
rect 43699 14241 43967 14249
tri 43967 14241 43975 14249 sw
tri 43699 14233 43707 14241 ne
rect 43707 14233 43975 14241
tri 43975 14233 43983 14241 sw
tri 43707 14225 43715 14233 ne
rect 43715 14225 43983 14233
tri 43983 14225 43991 14233 sw
tri 43715 14217 43723 14225 ne
rect 43723 14217 43991 14225
tri 43991 14217 43999 14225 sw
rect 70802 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43723 14209 43731 14217 ne
rect 43731 14209 43999 14217
tri 43999 14209 44007 14217 sw
tri 43731 14201 43739 14209 ne
rect 43739 14201 44007 14209
tri 44007 14201 44015 14209 sw
tri 43739 14193 43747 14201 ne
rect 43747 14200 44015 14201
rect 43747 14193 43878 14200
tri 43747 14185 43755 14193 ne
rect 43755 14185 43878 14193
tri 43755 14177 43763 14185 ne
rect 43763 14177 43878 14185
tri 43763 14169 43771 14177 ne
rect 43771 14169 43878 14177
tri 43771 14161 43779 14169 ne
rect 43779 14161 43878 14169
tri 43779 14153 43787 14161 ne
rect 43787 14154 43878 14161
rect 43924 14193 44015 14200
tri 44015 14193 44023 14201 sw
rect 43924 14185 44023 14193
tri 44023 14185 44031 14193 sw
rect 43924 14177 44031 14185
tri 44031 14177 44039 14185 sw
rect 43924 14169 44039 14177
tri 44039 14169 44047 14177 sw
rect 43924 14161 44047 14169
tri 44047 14161 44055 14169 sw
rect 70802 14164 71000 14222
rect 43924 14154 44055 14161
rect 43787 14153 44055 14154
tri 44055 14153 44063 14161 sw
tri 43787 14145 43795 14153 ne
rect 43795 14145 44063 14153
tri 44063 14145 44071 14153 sw
tri 43795 14137 43803 14145 ne
rect 43803 14141 44071 14145
tri 44071 14141 44075 14145 sw
rect 43803 14137 44075 14141
tri 43803 14130 43810 14137 ne
rect 43810 14133 44075 14137
tri 44075 14133 44083 14141 sw
rect 43810 14130 44083 14133
tri 43810 14122 43818 14130 ne
rect 43818 14125 44083 14130
tri 44083 14125 44091 14133 sw
rect 43818 14122 44091 14125
tri 43818 14114 43826 14122 ne
rect 43826 14117 44091 14122
tri 44091 14117 44099 14125 sw
rect 70802 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
rect 43826 14114 44099 14117
tri 43826 14106 43834 14114 ne
rect 43834 14109 44099 14114
tri 44099 14109 44107 14117 sw
rect 43834 14106 44107 14109
tri 43834 14098 43842 14106 ne
rect 43842 14101 44107 14106
tri 44107 14101 44115 14109 sw
rect 43842 14098 44115 14101
tri 43842 14090 43850 14098 ne
rect 43850 14093 44115 14098
tri 44115 14093 44123 14101 sw
rect 43850 14090 44123 14093
tri 43850 14082 43858 14090 ne
rect 43858 14085 44123 14090
tri 44123 14085 44131 14093 sw
rect 43858 14082 44131 14085
tri 43858 14074 43866 14082 ne
rect 43866 14077 44131 14082
tri 44131 14077 44139 14085 sw
rect 43866 14074 44139 14077
tri 43866 14066 43874 14074 ne
rect 43874 14069 44139 14074
tri 44139 14069 44147 14077 sw
rect 43874 14068 44147 14069
rect 43874 14066 44010 14068
tri 43874 14058 43882 14066 ne
rect 43882 14058 44010 14066
tri 43882 14050 43890 14058 ne
rect 43890 14050 44010 14058
tri 43890 14042 43898 14050 ne
rect 43898 14042 44010 14050
tri 43898 14034 43906 14042 ne
rect 43906 14034 44010 14042
tri 43906 14026 43914 14034 ne
rect 43914 14026 44010 14034
tri 43914 14018 43922 14026 ne
rect 43922 14022 44010 14026
rect 44056 14066 44147 14068
tri 44147 14066 44150 14069 sw
rect 44056 14058 44150 14066
tri 44150 14058 44158 14066 sw
rect 70802 14060 71000 14118
rect 44056 14050 44158 14058
tri 44158 14050 44166 14058 sw
rect 44056 14042 44166 14050
tri 44166 14042 44174 14050 sw
rect 44056 14034 44174 14042
tri 44174 14034 44182 14042 sw
rect 44056 14026 44182 14034
tri 44182 14026 44190 14034 sw
rect 44056 14022 44190 14026
rect 43922 14018 44190 14022
tri 44190 14018 44198 14026 sw
tri 43922 14010 43930 14018 ne
rect 43930 14010 44198 14018
tri 44198 14010 44206 14018 sw
rect 70802 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
tri 43930 14002 43938 14010 ne
rect 43938 14002 44206 14010
tri 44206 14002 44214 14010 sw
tri 43938 13994 43946 14002 ne
rect 43946 13994 44214 14002
tri 44214 13994 44222 14002 sw
tri 43946 13986 43954 13994 ne
rect 43954 13986 44222 13994
tri 44222 13986 44230 13994 sw
tri 43954 13978 43962 13986 ne
rect 43962 13978 44230 13986
tri 44230 13978 44238 13986 sw
tri 43962 13970 43970 13978 ne
rect 43970 13970 44238 13978
tri 44238 13970 44246 13978 sw
tri 43970 13962 43978 13970 ne
rect 43978 13962 44246 13970
tri 44246 13962 44254 13970 sw
tri 43978 13954 43986 13962 ne
rect 43986 13954 44254 13962
tri 44254 13954 44262 13962 sw
rect 70802 13956 71000 14014
tri 43986 13946 43994 13954 ne
rect 43994 13946 44262 13954
tri 44262 13946 44270 13954 sw
tri 43994 13938 44002 13946 ne
rect 44002 13938 44270 13946
tri 44270 13938 44278 13946 sw
tri 44002 13930 44010 13938 ne
rect 44010 13936 44278 13938
rect 44010 13930 44142 13936
tri 44010 13922 44018 13930 ne
rect 44018 13922 44142 13930
tri 44018 13914 44026 13922 ne
rect 44026 13914 44142 13922
tri 44026 13906 44034 13914 ne
rect 44034 13906 44142 13914
tri 44034 13898 44042 13906 ne
rect 44042 13898 44142 13906
tri 44042 13890 44050 13898 ne
rect 44050 13890 44142 13898
rect 44188 13930 44278 13936
tri 44278 13930 44286 13938 sw
rect 44188 13922 44286 13930
tri 44286 13922 44294 13930 sw
rect 44188 13914 44294 13922
tri 44294 13914 44302 13922 sw
rect 44188 13906 44302 13914
tri 44302 13906 44310 13914 sw
rect 70802 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 44188 13898 44310 13906
tri 44310 13898 44318 13906 sw
rect 44188 13890 44318 13898
tri 44318 13890 44326 13898 sw
tri 44050 13882 44058 13890 ne
rect 44058 13882 44326 13890
tri 44326 13882 44334 13890 sw
tri 44058 13874 44066 13882 ne
rect 44066 13874 44334 13882
tri 44334 13874 44342 13882 sw
tri 44066 13866 44074 13874 ne
rect 44074 13866 44342 13874
tri 44342 13866 44350 13874 sw
tri 44074 13862 44078 13866 ne
rect 44078 13862 44350 13866
tri 44078 13854 44086 13862 ne
rect 44086 13858 44350 13862
tri 44350 13858 44358 13866 sw
rect 44086 13854 44358 13858
tri 44086 13846 44094 13854 ne
rect 44094 13850 44358 13854
tri 44358 13850 44366 13858 sw
rect 70802 13852 71000 13910
rect 44094 13846 44366 13850
tri 44094 13838 44102 13846 ne
rect 44102 13842 44366 13846
tri 44366 13842 44374 13850 sw
rect 44102 13838 44374 13842
tri 44102 13830 44110 13838 ne
rect 44110 13834 44374 13838
tri 44374 13834 44382 13842 sw
rect 44110 13830 44382 13834
tri 44110 13822 44118 13830 ne
rect 44118 13826 44382 13830
tri 44382 13826 44390 13834 sw
rect 44118 13822 44390 13826
tri 44118 13814 44126 13822 ne
rect 44126 13818 44390 13822
tri 44390 13818 44398 13826 sw
rect 44126 13814 44398 13818
tri 44126 13806 44134 13814 ne
rect 44134 13811 44398 13814
tri 44398 13811 44405 13818 sw
rect 44134 13806 44405 13811
tri 44134 13798 44142 13806 ne
rect 44142 13804 44405 13806
rect 44142 13798 44274 13804
tri 44142 13795 44145 13798 ne
rect 44145 13795 44274 13798
tri 44145 13793 44147 13795 ne
rect 44147 13793 44274 13795
tri 44147 13787 44153 13793 ne
rect 44153 13787 44274 13793
tri 44153 13779 44161 13787 ne
rect 44161 13779 44274 13787
tri 44161 13771 44169 13779 ne
rect 44169 13771 44274 13779
tri 44169 13763 44177 13771 ne
rect 44177 13763 44274 13771
tri 44177 13755 44185 13763 ne
rect 44185 13758 44274 13763
rect 44320 13803 44405 13804
tri 44405 13803 44413 13811 sw
rect 70802 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 44320 13795 44413 13803
tri 44413 13795 44421 13803 sw
rect 44320 13787 44421 13795
tri 44421 13787 44429 13795 sw
rect 44320 13779 44429 13787
tri 44429 13779 44437 13787 sw
rect 44320 13771 44437 13779
tri 44437 13771 44445 13779 sw
rect 44320 13763 44445 13771
tri 44445 13763 44453 13771 sw
rect 44320 13758 44453 13763
rect 44185 13755 44453 13758
tri 44453 13755 44461 13763 sw
tri 44185 13747 44193 13755 ne
rect 44193 13747 44461 13755
tri 44461 13747 44469 13755 sw
rect 70802 13748 71000 13806
tri 44193 13739 44201 13747 ne
rect 44201 13739 44469 13747
tri 44469 13739 44477 13747 sw
tri 44201 13731 44209 13739 ne
rect 44209 13734 44477 13739
tri 44477 13734 44482 13739 sw
rect 44209 13731 44482 13734
tri 44209 13723 44217 13731 ne
rect 44217 13726 44482 13731
tri 44482 13726 44490 13734 sw
rect 44217 13723 44490 13726
tri 44217 13722 44218 13723 ne
rect 44218 13722 44490 13723
tri 44218 13714 44226 13722 ne
rect 44226 13718 44490 13722
tri 44490 13718 44498 13726 sw
rect 44226 13714 44498 13718
tri 44226 13706 44234 13714 ne
rect 44234 13710 44498 13714
tri 44498 13710 44506 13718 sw
rect 44234 13706 44506 13710
tri 44234 13698 44242 13706 ne
rect 44242 13702 44506 13706
tri 44506 13702 44514 13710 sw
rect 70802 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
rect 44242 13698 44514 13702
tri 44242 13690 44250 13698 ne
rect 44250 13694 44514 13698
tri 44514 13694 44522 13702 sw
rect 44250 13690 44522 13694
tri 44250 13682 44258 13690 ne
rect 44258 13686 44522 13690
tri 44522 13686 44530 13694 sw
rect 44258 13682 44530 13686
tri 44258 13674 44266 13682 ne
rect 44266 13678 44530 13682
tri 44530 13678 44538 13686 sw
rect 44266 13674 44538 13678
tri 44266 13666 44274 13674 ne
rect 44274 13672 44538 13674
rect 44274 13666 44406 13672
tri 44274 13658 44282 13666 ne
rect 44282 13658 44406 13666
tri 44282 13650 44290 13658 ne
rect 44290 13650 44406 13658
tri 44290 13642 44298 13650 ne
rect 44298 13642 44406 13650
tri 44298 13634 44306 13642 ne
rect 44306 13634 44406 13642
tri 44306 13626 44314 13634 ne
rect 44314 13626 44406 13634
rect 44452 13670 44538 13672
tri 44538 13670 44546 13678 sw
rect 44452 13662 44546 13670
tri 44546 13662 44554 13670 sw
rect 44452 13654 44554 13662
tri 44554 13654 44562 13662 sw
rect 44452 13646 44562 13654
tri 44562 13646 44570 13654 sw
rect 44452 13638 44570 13646
tri 44570 13638 44578 13646 sw
rect 70802 13644 71000 13702
rect 44452 13630 44578 13638
tri 44578 13630 44586 13638 sw
rect 44452 13626 44586 13630
tri 44314 13618 44322 13626 ne
rect 44322 13623 44586 13626
tri 44586 13623 44593 13630 sw
rect 44322 13618 44593 13623
tri 44322 13610 44330 13618 ne
rect 44330 13615 44593 13618
tri 44593 13615 44601 13623 sw
rect 44330 13610 44601 13615
tri 44330 13602 44338 13610 ne
rect 44338 13607 44601 13610
tri 44601 13607 44609 13615 sw
rect 44338 13602 44609 13607
tri 44338 13594 44346 13602 ne
rect 44346 13599 44609 13602
tri 44609 13599 44617 13607 sw
rect 44346 13594 44617 13599
tri 44346 13586 44354 13594 ne
rect 44354 13591 44617 13594
tri 44617 13591 44625 13599 sw
rect 70802 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44354 13586 44625 13591
tri 44354 13578 44362 13586 ne
rect 44362 13583 44625 13586
tri 44625 13583 44633 13591 sw
rect 44362 13578 44633 13583
tri 44362 13570 44370 13578 ne
rect 44370 13575 44633 13578
tri 44633 13575 44641 13583 sw
rect 44370 13570 44641 13575
tri 44370 13562 44378 13570 ne
rect 44378 13567 44641 13570
tri 44641 13567 44649 13575 sw
rect 44378 13562 44649 13567
tri 44378 13554 44386 13562 ne
rect 44386 13559 44649 13562
tri 44649 13559 44657 13567 sw
rect 44386 13554 44657 13559
tri 44386 13546 44394 13554 ne
rect 44394 13551 44657 13554
tri 44657 13551 44665 13559 sw
rect 44394 13546 44665 13551
tri 44394 13538 44402 13546 ne
rect 44402 13543 44665 13546
tri 44665 13543 44673 13551 sw
rect 44402 13540 44673 13543
rect 44402 13538 44538 13540
tri 44402 13534 44406 13538 ne
rect 44406 13534 44538 13538
tri 44406 13530 44410 13534 ne
rect 44410 13530 44538 13534
tri 44410 13522 44418 13530 ne
rect 44418 13522 44538 13530
tri 44418 13514 44426 13522 ne
rect 44426 13514 44538 13522
tri 44426 13506 44434 13514 ne
rect 44434 13506 44538 13514
tri 44434 13498 44442 13506 ne
rect 44442 13498 44538 13506
tri 44442 13490 44450 13498 ne
rect 44450 13494 44538 13498
rect 44584 13535 44673 13540
tri 44673 13535 44681 13543 sw
rect 70802 13540 71000 13598
rect 44584 13527 44681 13535
tri 44681 13527 44689 13535 sw
rect 44584 13519 44689 13527
tri 44689 13519 44697 13527 sw
rect 44584 13511 44697 13519
tri 44697 13511 44705 13519 sw
rect 44584 13503 44705 13511
tri 44705 13503 44713 13511 sw
rect 44584 13495 44713 13503
tri 44713 13495 44721 13503 sw
rect 44584 13494 44721 13495
rect 44450 13490 44721 13494
tri 44450 13482 44458 13490 ne
rect 44458 13487 44721 13490
tri 44721 13487 44729 13495 sw
rect 70802 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
rect 44458 13482 44729 13487
tri 44458 13474 44466 13482 ne
rect 44466 13479 44729 13482
tri 44729 13479 44737 13487 sw
rect 44466 13474 44737 13479
tri 44466 13466 44474 13474 ne
rect 44474 13471 44737 13474
tri 44737 13471 44745 13479 sw
rect 44474 13466 44745 13471
tri 44474 13458 44482 13466 ne
rect 44482 13463 44745 13466
tri 44745 13463 44753 13471 sw
rect 44482 13458 44753 13463
tri 44482 13450 44490 13458 ne
rect 44490 13455 44753 13458
tri 44753 13455 44761 13463 sw
rect 44490 13450 44761 13455
tri 44490 13442 44498 13450 ne
rect 44498 13447 44761 13450
tri 44761 13447 44769 13455 sw
rect 44498 13442 44769 13447
tri 44498 13434 44506 13442 ne
rect 44506 13439 44769 13442
tri 44769 13439 44777 13447 sw
rect 44506 13434 44777 13439
tri 44506 13426 44514 13434 ne
rect 44514 13431 44777 13434
tri 44777 13431 44785 13439 sw
rect 70802 13436 71000 13494
rect 44514 13426 44785 13431
tri 44514 13418 44522 13426 ne
rect 44522 13423 44785 13426
tri 44785 13423 44793 13431 sw
rect 44522 13418 44793 13423
tri 44522 13410 44530 13418 ne
rect 44530 13415 44793 13418
tri 44793 13415 44801 13423 sw
rect 44530 13410 44801 13415
tri 44530 13403 44537 13410 ne
rect 44537 13408 44801 13410
rect 44537 13403 44670 13408
tri 44537 13395 44545 13403 ne
rect 44545 13395 44670 13403
tri 44545 13387 44553 13395 ne
rect 44553 13387 44670 13395
tri 44553 13379 44561 13387 ne
rect 44561 13379 44670 13387
tri 44561 13371 44569 13379 ne
rect 44569 13371 44670 13379
tri 44569 13363 44577 13371 ne
rect 44577 13363 44670 13371
tri 44577 13355 44585 13363 ne
rect 44585 13362 44670 13363
rect 44716 13407 44801 13408
tri 44801 13407 44809 13415 sw
rect 44716 13399 44809 13407
tri 44809 13399 44817 13407 sw
rect 44716 13391 44817 13399
tri 44817 13391 44825 13399 sw
rect 44716 13383 44825 13391
tri 44825 13383 44833 13391 sw
rect 70802 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13375 44833 13383
tri 44833 13375 44841 13383 sw
rect 44716 13367 44841 13375
tri 44841 13367 44849 13375 sw
rect 44716 13362 44849 13367
rect 44585 13359 44849 13362
tri 44849 13359 44857 13367 sw
rect 44585 13355 44857 13359
tri 44585 13347 44593 13355 ne
rect 44593 13351 44857 13355
tri 44857 13351 44865 13359 sw
rect 44593 13347 44865 13351
tri 44593 13339 44601 13347 ne
rect 44601 13343 44865 13347
tri 44865 13343 44873 13351 sw
rect 44601 13339 44873 13343
tri 44601 13331 44609 13339 ne
rect 44609 13335 44873 13339
tri 44873 13335 44881 13343 sw
rect 44609 13331 44881 13335
tri 44609 13323 44617 13331 ne
rect 44617 13327 44881 13331
tri 44881 13327 44889 13335 sw
rect 44617 13323 44889 13327
tri 44617 13315 44625 13323 ne
rect 44625 13319 44889 13323
tri 44889 13319 44897 13327 sw
rect 44625 13315 44897 13319
tri 44625 13307 44633 13315 ne
rect 44633 13311 44897 13315
tri 44897 13311 44905 13319 sw
rect 44633 13307 44905 13311
tri 44633 13299 44641 13307 ne
rect 44641 13303 44905 13307
tri 44905 13303 44913 13311 sw
rect 44641 13299 44913 13303
tri 44641 13291 44649 13299 ne
rect 44649 13295 44913 13299
tri 44913 13295 44921 13303 sw
rect 44649 13291 44921 13295
tri 44921 13291 44925 13295 sw
rect 70802 13291 71000 13390
tri 44649 13283 44657 13291 ne
rect 44657 13283 71000 13291
tri 44657 13275 44665 13283 ne
rect 44665 13275 71000 13283
tri 44665 13267 44673 13275 ne
rect 44673 13269 71000 13275
rect 44673 13267 45088 13269
tri 44673 13259 44681 13267 ne
rect 44681 13259 45088 13267
tri 44681 13251 44689 13259 ne
rect 44689 13256 45088 13259
rect 44689 13251 44850 13256
tri 44689 13243 44697 13251 ne
rect 44697 13243 44850 13251
tri 44697 13235 44705 13243 ne
rect 44705 13235 44850 13243
tri 44705 13227 44713 13235 ne
rect 44713 13227 44850 13235
tri 44713 13219 44721 13227 ne
rect 44721 13219 44850 13227
tri 44721 13211 44729 13219 ne
rect 44729 13211 44850 13219
tri 44729 13203 44737 13211 ne
rect 44737 13210 44850 13211
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44737 13203 71000 13210
tri 44737 13195 44745 13203 ne
rect 44745 13195 71000 13203
tri 44745 13187 44753 13195 ne
rect 44753 13187 71000 13195
tri 44753 13181 44759 13187 ne
rect 44759 13181 71000 13187
tri 44759 13173 44767 13181 ne
rect 44767 13173 71000 13181
tri 44767 13165 44775 13173 ne
rect 44775 13165 71000 13173
tri 44775 13157 44783 13165 ne
rect 44783 13157 45088 13165
tri 44783 13149 44791 13157 ne
rect 44791 13149 45088 13157
tri 44791 13141 44799 13149 ne
rect 44799 13141 45088 13149
tri 44799 13133 44807 13141 ne
rect 44807 13133 45088 13141
tri 44807 13125 44815 13133 ne
rect 44815 13125 45088 13133
tri 44815 13117 44823 13125 ne
rect 44823 13119 45088 13125
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44823 13117 71000 13119
tri 44823 13109 44831 13117 ne
rect 44831 13109 71000 13117
tri 44831 13101 44839 13109 ne
rect 44839 13101 71000 13109
tri 44839 13097 44843 13101 ne
rect 44843 13097 71000 13101
<< psubdiffcont >>
rect 13119 70929 13165 70975
rect 13223 70929 13269 70975
rect 13377 70929 13423 70975
rect 13481 70929 13527 70975
rect 13585 70929 13631 70975
rect 13689 70929 13735 70975
rect 13793 70929 13839 70975
rect 13897 70929 13943 70975
rect 14001 70929 14047 70975
rect 14105 70929 14151 70975
rect 14209 70929 14255 70975
rect 14313 70929 14359 70975
rect 14417 70929 14463 70975
rect 14521 70929 14567 70975
rect 14625 70929 14671 70975
rect 14729 70929 14775 70975
rect 14833 70929 14879 70975
rect 14937 70929 14983 70975
rect 15041 70929 15087 70975
rect 15145 70929 15191 70975
rect 15249 70929 15295 70975
rect 15353 70929 15399 70975
rect 15457 70929 15503 70975
rect 15561 70929 15607 70975
rect 15665 70929 15711 70975
rect 15769 70929 15815 70975
rect 15873 70929 15919 70975
rect 15977 70929 16023 70975
rect 16081 70929 16127 70975
rect 16185 70929 16231 70975
rect 16289 70929 16335 70975
rect 16393 70929 16439 70975
rect 16497 70929 16543 70975
rect 16601 70929 16647 70975
rect 16705 70929 16751 70975
rect 16809 70929 16855 70975
rect 16913 70929 16959 70975
rect 17017 70929 17063 70975
rect 17121 70929 17167 70975
rect 17225 70929 17271 70975
rect 17329 70929 17375 70975
rect 17433 70929 17479 70975
rect 17537 70929 17583 70975
rect 17641 70929 17687 70975
rect 17745 70929 17791 70975
rect 17849 70929 17895 70975
rect 17953 70929 17999 70975
rect 18057 70929 18103 70975
rect 18161 70929 18207 70975
rect 18265 70929 18311 70975
rect 18369 70929 18415 70975
rect 18473 70929 18519 70975
rect 18577 70929 18623 70975
rect 18681 70929 18727 70975
rect 18785 70929 18831 70975
rect 18889 70929 18935 70975
rect 18993 70929 19039 70975
rect 19097 70929 19143 70975
rect 19201 70929 19247 70975
rect 19305 70929 19351 70975
rect 19409 70929 19455 70975
rect 19513 70929 19559 70975
rect 19617 70929 19663 70975
rect 19721 70929 19767 70975
rect 19825 70929 19871 70975
rect 19929 70929 19975 70975
rect 20033 70929 20079 70975
rect 20137 70929 20183 70975
rect 20241 70929 20287 70975
rect 20345 70929 20391 70975
rect 20449 70929 20495 70975
rect 20553 70929 20599 70975
rect 20657 70929 20703 70975
rect 20761 70929 20807 70975
rect 20865 70929 20911 70975
rect 20969 70929 21015 70975
rect 21073 70929 21119 70975
rect 21177 70929 21223 70975
rect 21281 70929 21327 70975
rect 21385 70929 21431 70975
rect 21489 70929 21535 70975
rect 21593 70929 21639 70975
rect 21697 70929 21743 70975
rect 21801 70929 21847 70975
rect 21905 70929 21951 70975
rect 22009 70929 22055 70975
rect 22113 70929 22159 70975
rect 22217 70929 22263 70975
rect 22321 70929 22367 70975
rect 22425 70929 22471 70975
rect 22529 70929 22575 70975
rect 22633 70929 22679 70975
rect 22737 70929 22783 70975
rect 22841 70929 22887 70975
rect 22945 70929 22991 70975
rect 23049 70929 23095 70975
rect 23153 70929 23199 70975
rect 23257 70929 23303 70975
rect 23361 70929 23407 70975
rect 23465 70929 23511 70975
rect 23569 70929 23615 70975
rect 23673 70929 23719 70975
rect 23777 70929 23823 70975
rect 23881 70929 23927 70975
rect 23985 70929 24031 70975
rect 24089 70929 24135 70975
rect 24193 70929 24239 70975
rect 24297 70929 24343 70975
rect 24401 70929 24447 70975
rect 24505 70929 24551 70975
rect 24609 70929 24655 70975
rect 24713 70929 24759 70975
rect 24817 70929 24863 70975
rect 24921 70929 24967 70975
rect 25025 70929 25071 70975
rect 25129 70929 25175 70975
rect 25233 70929 25279 70975
rect 25337 70929 25383 70975
rect 25441 70929 25487 70975
rect 25545 70929 25591 70975
rect 25649 70929 25695 70975
rect 25753 70929 25799 70975
rect 25857 70929 25903 70975
rect 25961 70929 26007 70975
rect 26065 70929 26111 70975
rect 26169 70929 26215 70975
rect 26273 70929 26319 70975
rect 26377 70929 26423 70975
rect 26481 70929 26527 70975
rect 26585 70929 26631 70975
rect 26689 70929 26735 70975
rect 26793 70929 26839 70975
rect 26897 70929 26943 70975
rect 27001 70929 27047 70975
rect 27105 70929 27151 70975
rect 27209 70929 27255 70975
rect 27313 70929 27359 70975
rect 27417 70929 27463 70975
rect 27521 70929 27567 70975
rect 27625 70929 27671 70975
rect 27729 70929 27775 70975
rect 27833 70929 27879 70975
rect 27937 70929 27983 70975
rect 28041 70929 28087 70975
rect 28145 70929 28191 70975
rect 28249 70929 28295 70975
rect 28353 70929 28399 70975
rect 28457 70929 28503 70975
rect 28561 70929 28607 70975
rect 28665 70929 28711 70975
rect 28769 70929 28815 70975
rect 28873 70929 28919 70975
rect 28977 70929 29023 70975
rect 29081 70929 29127 70975
rect 29185 70929 29231 70975
rect 29289 70929 29335 70975
rect 29393 70929 29439 70975
rect 29497 70929 29543 70975
rect 29601 70929 29647 70975
rect 29705 70929 29751 70975
rect 29809 70929 29855 70975
rect 29913 70929 29959 70975
rect 30017 70929 30063 70975
rect 30121 70929 30167 70975
rect 30225 70929 30271 70975
rect 30329 70929 30375 70975
rect 30433 70929 30479 70975
rect 30537 70929 30583 70975
rect 30641 70929 30687 70975
rect 30745 70929 30791 70975
rect 30849 70929 30895 70975
rect 30953 70929 30999 70975
rect 31057 70929 31103 70975
rect 31161 70929 31207 70975
rect 31265 70929 31311 70975
rect 31369 70929 31415 70975
rect 31473 70929 31519 70975
rect 31577 70929 31623 70975
rect 31681 70929 31727 70975
rect 31785 70929 31831 70975
rect 31889 70929 31935 70975
rect 31993 70929 32039 70975
rect 32097 70929 32143 70975
rect 32201 70929 32247 70975
rect 32305 70929 32351 70975
rect 32409 70929 32455 70975
rect 32513 70929 32559 70975
rect 32617 70929 32663 70975
rect 32721 70929 32767 70975
rect 32825 70929 32871 70975
rect 32929 70929 32975 70975
rect 33033 70929 33079 70975
rect 33137 70929 33183 70975
rect 33241 70929 33287 70975
rect 33345 70929 33391 70975
rect 33449 70929 33495 70975
rect 33553 70929 33599 70975
rect 33657 70929 33703 70975
rect 33761 70929 33807 70975
rect 33865 70929 33911 70975
rect 33969 70929 34015 70975
rect 34073 70929 34119 70975
rect 34177 70929 34223 70975
rect 34281 70929 34327 70975
rect 34385 70929 34431 70975
rect 34489 70929 34535 70975
rect 34593 70929 34639 70975
rect 34697 70929 34743 70975
rect 34801 70929 34847 70975
rect 34905 70929 34951 70975
rect 35009 70929 35055 70975
rect 35113 70929 35159 70975
rect 35217 70929 35263 70975
rect 35321 70929 35367 70975
rect 35425 70929 35471 70975
rect 35529 70929 35575 70975
rect 35633 70929 35679 70975
rect 35737 70929 35783 70975
rect 35841 70929 35887 70975
rect 35945 70929 35991 70975
rect 36049 70929 36095 70975
rect 36153 70929 36199 70975
rect 36257 70929 36303 70975
rect 36361 70929 36407 70975
rect 36465 70929 36511 70975
rect 36569 70929 36615 70975
rect 36673 70929 36719 70975
rect 36777 70929 36823 70975
rect 36881 70929 36927 70975
rect 36985 70929 37031 70975
rect 37089 70929 37135 70975
rect 37193 70929 37239 70975
rect 37297 70929 37343 70975
rect 37401 70929 37447 70975
rect 37505 70929 37551 70975
rect 37609 70929 37655 70975
rect 37713 70929 37759 70975
rect 37817 70929 37863 70975
rect 37921 70929 37967 70975
rect 38025 70929 38071 70975
rect 38129 70929 38175 70975
rect 38233 70929 38279 70975
rect 38337 70929 38383 70975
rect 38441 70929 38487 70975
rect 38545 70929 38591 70975
rect 38649 70929 38695 70975
rect 38753 70929 38799 70975
rect 38857 70929 38903 70975
rect 38961 70929 39007 70975
rect 39065 70929 39111 70975
rect 39169 70929 39215 70975
rect 39273 70929 39319 70975
rect 39377 70929 39423 70975
rect 39481 70929 39527 70975
rect 39585 70929 39631 70975
rect 39689 70929 39735 70975
rect 39793 70929 39839 70975
rect 39897 70929 39943 70975
rect 40001 70929 40047 70975
rect 40105 70929 40151 70975
rect 40209 70929 40255 70975
rect 40313 70929 40359 70975
rect 40417 70929 40463 70975
rect 40521 70929 40567 70975
rect 40625 70929 40671 70975
rect 40729 70929 40775 70975
rect 40833 70929 40879 70975
rect 40937 70929 40983 70975
rect 41041 70929 41087 70975
rect 41145 70929 41191 70975
rect 41249 70929 41295 70975
rect 41353 70929 41399 70975
rect 41457 70929 41503 70975
rect 41561 70929 41607 70975
rect 41665 70929 41711 70975
rect 41769 70929 41815 70975
rect 41873 70929 41919 70975
rect 41977 70929 42023 70975
rect 42081 70929 42127 70975
rect 42185 70929 42231 70975
rect 42289 70929 42335 70975
rect 42393 70929 42439 70975
rect 42497 70929 42543 70975
rect 42601 70929 42647 70975
rect 42705 70929 42751 70975
rect 42809 70929 42855 70975
rect 42913 70929 42959 70975
rect 43017 70929 43063 70975
rect 43121 70929 43167 70975
rect 43225 70929 43271 70975
rect 43329 70929 43375 70975
rect 43433 70929 43479 70975
rect 43537 70929 43583 70975
rect 43641 70929 43687 70975
rect 43745 70929 43791 70975
rect 43849 70929 43895 70975
rect 43953 70929 43999 70975
rect 44057 70929 44103 70975
rect 44161 70929 44207 70975
rect 44265 70929 44311 70975
rect 44369 70929 44415 70975
rect 44473 70929 44519 70975
rect 44577 70929 44623 70975
rect 44681 70929 44727 70975
rect 44785 70929 44831 70975
rect 44889 70929 44935 70975
rect 44993 70929 45039 70975
rect 45097 70929 45143 70975
rect 45201 70929 45247 70975
rect 45305 70929 45351 70975
rect 45409 70929 45455 70975
rect 45513 70929 45559 70975
rect 45617 70929 45663 70975
rect 45721 70929 45767 70975
rect 45825 70929 45871 70975
rect 45929 70929 45975 70975
rect 46033 70929 46079 70975
rect 46137 70929 46183 70975
rect 46241 70929 46287 70975
rect 46345 70929 46391 70975
rect 46449 70929 46495 70975
rect 46553 70929 46599 70975
rect 46657 70929 46703 70975
rect 46761 70929 46807 70975
rect 46865 70929 46911 70975
rect 46969 70929 47015 70975
rect 47073 70929 47119 70975
rect 47177 70929 47223 70975
rect 47281 70929 47327 70975
rect 47385 70929 47431 70975
rect 47489 70929 47535 70975
rect 47593 70929 47639 70975
rect 47697 70929 47743 70975
rect 47801 70929 47847 70975
rect 47905 70929 47951 70975
rect 48009 70929 48055 70975
rect 48113 70929 48159 70975
rect 48217 70929 48263 70975
rect 48321 70929 48367 70975
rect 48425 70929 48471 70975
rect 48529 70929 48575 70975
rect 48633 70929 48679 70975
rect 48737 70929 48783 70975
rect 48841 70929 48887 70975
rect 48945 70929 48991 70975
rect 49049 70929 49095 70975
rect 49153 70929 49199 70975
rect 49257 70929 49303 70975
rect 49361 70929 49407 70975
rect 49465 70929 49511 70975
rect 49569 70929 49615 70975
rect 49673 70929 49719 70975
rect 49777 70929 49823 70975
rect 49881 70929 49927 70975
rect 49985 70929 50031 70975
rect 50089 70929 50135 70975
rect 50193 70929 50239 70975
rect 50297 70929 50343 70975
rect 50401 70929 50447 70975
rect 50505 70929 50551 70975
rect 50609 70929 50655 70975
rect 50713 70929 50759 70975
rect 50817 70929 50863 70975
rect 50921 70929 50967 70975
rect 51025 70929 51071 70975
rect 51129 70929 51175 70975
rect 51233 70929 51279 70975
rect 51337 70929 51383 70975
rect 51441 70929 51487 70975
rect 51545 70929 51591 70975
rect 51649 70929 51695 70975
rect 51753 70929 51799 70975
rect 51857 70929 51903 70975
rect 51961 70929 52007 70975
rect 52065 70929 52111 70975
rect 52169 70929 52215 70975
rect 52273 70929 52319 70975
rect 52377 70929 52423 70975
rect 52481 70929 52527 70975
rect 52585 70929 52631 70975
rect 52689 70929 52735 70975
rect 52793 70929 52839 70975
rect 52897 70929 52943 70975
rect 53001 70929 53047 70975
rect 53105 70929 53151 70975
rect 53209 70929 53255 70975
rect 53313 70929 53359 70975
rect 53417 70929 53463 70975
rect 53521 70929 53567 70975
rect 53625 70929 53671 70975
rect 53729 70929 53775 70975
rect 53833 70929 53879 70975
rect 53937 70929 53983 70975
rect 54041 70929 54087 70975
rect 54145 70929 54191 70975
rect 54249 70929 54295 70975
rect 54353 70929 54399 70975
rect 54457 70929 54503 70975
rect 54561 70929 54607 70975
rect 54665 70929 54711 70975
rect 54769 70929 54815 70975
rect 54873 70929 54919 70975
rect 54977 70929 55023 70975
rect 55081 70929 55127 70975
rect 55185 70929 55231 70975
rect 55289 70929 55335 70975
rect 55393 70929 55439 70975
rect 55497 70929 55543 70975
rect 55601 70929 55647 70975
rect 55705 70929 55751 70975
rect 55809 70929 55855 70975
rect 55913 70929 55959 70975
rect 56017 70929 56063 70975
rect 56121 70929 56167 70975
rect 56225 70929 56271 70975
rect 56329 70929 56375 70975
rect 56433 70929 56479 70975
rect 56537 70929 56583 70975
rect 56641 70929 56687 70975
rect 56745 70929 56791 70975
rect 56849 70929 56895 70975
rect 56953 70929 56999 70975
rect 57057 70929 57103 70975
rect 57161 70929 57207 70975
rect 57265 70929 57311 70975
rect 57369 70929 57415 70975
rect 57473 70929 57519 70975
rect 57577 70929 57623 70975
rect 57681 70929 57727 70975
rect 57785 70929 57831 70975
rect 57889 70929 57935 70975
rect 57993 70929 58039 70975
rect 58097 70929 58143 70975
rect 58201 70929 58247 70975
rect 58305 70929 58351 70975
rect 58409 70929 58455 70975
rect 58513 70929 58559 70975
rect 58617 70929 58663 70975
rect 58721 70929 58767 70975
rect 58825 70929 58871 70975
rect 58929 70929 58975 70975
rect 59033 70929 59079 70975
rect 59137 70929 59183 70975
rect 59241 70929 59287 70975
rect 59345 70929 59391 70975
rect 59449 70929 59495 70975
rect 59553 70929 59599 70975
rect 59657 70929 59703 70975
rect 59761 70929 59807 70975
rect 59865 70929 59911 70975
rect 59969 70929 60015 70975
rect 60073 70929 60119 70975
rect 60177 70929 60223 70975
rect 60281 70929 60327 70975
rect 60385 70929 60431 70975
rect 60489 70929 60535 70975
rect 60593 70929 60639 70975
rect 60697 70929 60743 70975
rect 60801 70929 60847 70975
rect 60905 70929 60951 70975
rect 61009 70929 61055 70975
rect 61113 70929 61159 70975
rect 61217 70929 61263 70975
rect 61321 70929 61367 70975
rect 61425 70929 61471 70975
rect 61529 70929 61575 70975
rect 61633 70929 61679 70975
rect 61737 70929 61783 70975
rect 61841 70929 61887 70975
rect 61945 70929 61991 70975
rect 62049 70929 62095 70975
rect 62153 70929 62199 70975
rect 62257 70929 62303 70975
rect 62361 70929 62407 70975
rect 62465 70929 62511 70975
rect 62569 70929 62615 70975
rect 62673 70929 62719 70975
rect 62777 70929 62823 70975
rect 62881 70929 62927 70975
rect 62985 70929 63031 70975
rect 63089 70929 63135 70975
rect 63193 70929 63239 70975
rect 63297 70929 63343 70975
rect 63401 70929 63447 70975
rect 63505 70929 63551 70975
rect 63609 70929 63655 70975
rect 63713 70929 63759 70975
rect 63817 70929 63863 70975
rect 63921 70929 63967 70975
rect 64025 70929 64071 70975
rect 64129 70929 64175 70975
rect 64233 70929 64279 70975
rect 64337 70929 64383 70975
rect 64441 70929 64487 70975
rect 64545 70929 64591 70975
rect 64649 70929 64695 70975
rect 64753 70929 64799 70975
rect 64857 70929 64903 70975
rect 64961 70929 65007 70975
rect 65065 70929 65111 70975
rect 65169 70929 65215 70975
rect 65273 70929 65319 70975
rect 65377 70929 65423 70975
rect 65481 70929 65527 70975
rect 65585 70929 65631 70975
rect 65689 70929 65735 70975
rect 65793 70929 65839 70975
rect 65897 70929 65943 70975
rect 66001 70929 66047 70975
rect 66105 70929 66151 70975
rect 66209 70929 66255 70975
rect 66313 70929 66359 70975
rect 66417 70929 66463 70975
rect 66521 70929 66567 70975
rect 66625 70929 66671 70975
rect 66729 70929 66775 70975
rect 66833 70929 66879 70975
rect 66937 70929 66983 70975
rect 67041 70929 67087 70975
rect 67145 70929 67191 70975
rect 67249 70929 67295 70975
rect 67353 70929 67399 70975
rect 67457 70929 67503 70975
rect 67561 70929 67607 70975
rect 67665 70929 67711 70975
rect 67769 70929 67815 70975
rect 67873 70929 67919 70975
rect 67977 70929 68023 70975
rect 68081 70929 68127 70975
rect 68185 70929 68231 70975
rect 68289 70929 68335 70975
rect 68393 70929 68439 70975
rect 68497 70929 68543 70975
rect 68601 70929 68647 70975
rect 68705 70929 68751 70975
rect 68809 70929 68855 70975
rect 68913 70929 68959 70975
rect 69017 70929 69063 70975
rect 69121 70929 69167 70975
rect 69225 70929 69271 70975
rect 69329 70929 69375 70975
rect 69433 70929 69479 70975
rect 69537 70929 69583 70975
rect 69641 70929 69687 70975
rect 69745 70929 69791 70975
rect 69849 70929 69895 70975
rect 13119 70825 13165 70871
rect 13223 70825 13269 70871
rect 13377 70825 13423 70871
rect 13481 70825 13527 70871
rect 13585 70825 13631 70871
rect 13689 70825 13735 70871
rect 13793 70825 13839 70871
rect 13897 70825 13943 70871
rect 14001 70825 14047 70871
rect 14105 70825 14151 70871
rect 14209 70825 14255 70871
rect 14313 70825 14359 70871
rect 14417 70825 14463 70871
rect 14521 70825 14567 70871
rect 14625 70825 14671 70871
rect 14729 70825 14775 70871
rect 14833 70825 14879 70871
rect 14937 70825 14983 70871
rect 15041 70825 15087 70871
rect 15145 70825 15191 70871
rect 15249 70825 15295 70871
rect 15353 70825 15399 70871
rect 15457 70825 15503 70871
rect 15561 70825 15607 70871
rect 15665 70825 15711 70871
rect 15769 70825 15815 70871
rect 15873 70825 15919 70871
rect 15977 70825 16023 70871
rect 16081 70825 16127 70871
rect 16185 70825 16231 70871
rect 16289 70825 16335 70871
rect 16393 70825 16439 70871
rect 16497 70825 16543 70871
rect 16601 70825 16647 70871
rect 16705 70825 16751 70871
rect 16809 70825 16855 70871
rect 16913 70825 16959 70871
rect 17017 70825 17063 70871
rect 17121 70825 17167 70871
rect 17225 70825 17271 70871
rect 17329 70825 17375 70871
rect 17433 70825 17479 70871
rect 17537 70825 17583 70871
rect 17641 70825 17687 70871
rect 17745 70825 17791 70871
rect 17849 70825 17895 70871
rect 17953 70825 17999 70871
rect 18057 70825 18103 70871
rect 18161 70825 18207 70871
rect 18265 70825 18311 70871
rect 18369 70825 18415 70871
rect 18473 70825 18519 70871
rect 18577 70825 18623 70871
rect 18681 70825 18727 70871
rect 18785 70825 18831 70871
rect 18889 70825 18935 70871
rect 18993 70825 19039 70871
rect 19097 70825 19143 70871
rect 19201 70825 19247 70871
rect 19305 70825 19351 70871
rect 19409 70825 19455 70871
rect 19513 70825 19559 70871
rect 19617 70825 19663 70871
rect 19721 70825 19767 70871
rect 19825 70825 19871 70871
rect 19929 70825 19975 70871
rect 20033 70825 20079 70871
rect 20137 70825 20183 70871
rect 20241 70825 20287 70871
rect 20345 70825 20391 70871
rect 20449 70825 20495 70871
rect 20553 70825 20599 70871
rect 20657 70825 20703 70871
rect 20761 70825 20807 70871
rect 20865 70825 20911 70871
rect 20969 70825 21015 70871
rect 21073 70825 21119 70871
rect 21177 70825 21223 70871
rect 21281 70825 21327 70871
rect 21385 70825 21431 70871
rect 21489 70825 21535 70871
rect 21593 70825 21639 70871
rect 21697 70825 21743 70871
rect 21801 70825 21847 70871
rect 21905 70825 21951 70871
rect 22009 70825 22055 70871
rect 22113 70825 22159 70871
rect 22217 70825 22263 70871
rect 22321 70825 22367 70871
rect 22425 70825 22471 70871
rect 22529 70825 22575 70871
rect 22633 70825 22679 70871
rect 22737 70825 22783 70871
rect 22841 70825 22887 70871
rect 22945 70825 22991 70871
rect 23049 70825 23095 70871
rect 23153 70825 23199 70871
rect 23257 70825 23303 70871
rect 23361 70825 23407 70871
rect 23465 70825 23511 70871
rect 23569 70825 23615 70871
rect 23673 70825 23719 70871
rect 23777 70825 23823 70871
rect 23881 70825 23927 70871
rect 23985 70825 24031 70871
rect 24089 70825 24135 70871
rect 24193 70825 24239 70871
rect 24297 70825 24343 70871
rect 24401 70825 24447 70871
rect 24505 70825 24551 70871
rect 24609 70825 24655 70871
rect 24713 70825 24759 70871
rect 24817 70825 24863 70871
rect 24921 70825 24967 70871
rect 25025 70825 25071 70871
rect 25129 70825 25175 70871
rect 25233 70825 25279 70871
rect 25337 70825 25383 70871
rect 25441 70825 25487 70871
rect 25545 70825 25591 70871
rect 25649 70825 25695 70871
rect 25753 70825 25799 70871
rect 25857 70825 25903 70871
rect 25961 70825 26007 70871
rect 26065 70825 26111 70871
rect 26169 70825 26215 70871
rect 26273 70825 26319 70871
rect 26377 70825 26423 70871
rect 26481 70825 26527 70871
rect 26585 70825 26631 70871
rect 26689 70825 26735 70871
rect 26793 70825 26839 70871
rect 26897 70825 26943 70871
rect 27001 70825 27047 70871
rect 27105 70825 27151 70871
rect 27209 70825 27255 70871
rect 27313 70825 27359 70871
rect 27417 70825 27463 70871
rect 27521 70825 27567 70871
rect 27625 70825 27671 70871
rect 27729 70825 27775 70871
rect 27833 70825 27879 70871
rect 27937 70825 27983 70871
rect 28041 70825 28087 70871
rect 28145 70825 28191 70871
rect 28249 70825 28295 70871
rect 28353 70825 28399 70871
rect 28457 70825 28503 70871
rect 28561 70825 28607 70871
rect 28665 70825 28711 70871
rect 28769 70825 28815 70871
rect 28873 70825 28919 70871
rect 28977 70825 29023 70871
rect 29081 70825 29127 70871
rect 29185 70825 29231 70871
rect 29289 70825 29335 70871
rect 29393 70825 29439 70871
rect 29497 70825 29543 70871
rect 29601 70825 29647 70871
rect 29705 70825 29751 70871
rect 29809 70825 29855 70871
rect 29913 70825 29959 70871
rect 30017 70825 30063 70871
rect 30121 70825 30167 70871
rect 30225 70825 30271 70871
rect 30329 70825 30375 70871
rect 30433 70825 30479 70871
rect 30537 70825 30583 70871
rect 30641 70825 30687 70871
rect 30745 70825 30791 70871
rect 30849 70825 30895 70871
rect 30953 70825 30999 70871
rect 31057 70825 31103 70871
rect 31161 70825 31207 70871
rect 31265 70825 31311 70871
rect 31369 70825 31415 70871
rect 31473 70825 31519 70871
rect 31577 70825 31623 70871
rect 31681 70825 31727 70871
rect 31785 70825 31831 70871
rect 31889 70825 31935 70871
rect 31993 70825 32039 70871
rect 32097 70825 32143 70871
rect 32201 70825 32247 70871
rect 32305 70825 32351 70871
rect 32409 70825 32455 70871
rect 32513 70825 32559 70871
rect 32617 70825 32663 70871
rect 32721 70825 32767 70871
rect 32825 70825 32871 70871
rect 32929 70825 32975 70871
rect 33033 70825 33079 70871
rect 33137 70825 33183 70871
rect 33241 70825 33287 70871
rect 33345 70825 33391 70871
rect 33449 70825 33495 70871
rect 33553 70825 33599 70871
rect 33657 70825 33703 70871
rect 33761 70825 33807 70871
rect 33865 70825 33911 70871
rect 33969 70825 34015 70871
rect 34073 70825 34119 70871
rect 34177 70825 34223 70871
rect 34281 70825 34327 70871
rect 34385 70825 34431 70871
rect 34489 70825 34535 70871
rect 34593 70825 34639 70871
rect 34697 70825 34743 70871
rect 34801 70825 34847 70871
rect 34905 70825 34951 70871
rect 35009 70825 35055 70871
rect 35113 70825 35159 70871
rect 35217 70825 35263 70871
rect 35321 70825 35367 70871
rect 35425 70825 35471 70871
rect 35529 70825 35575 70871
rect 35633 70825 35679 70871
rect 35737 70825 35783 70871
rect 35841 70825 35887 70871
rect 35945 70825 35991 70871
rect 36049 70825 36095 70871
rect 36153 70825 36199 70871
rect 36257 70825 36303 70871
rect 36361 70825 36407 70871
rect 36465 70825 36511 70871
rect 36569 70825 36615 70871
rect 36673 70825 36719 70871
rect 36777 70825 36823 70871
rect 36881 70825 36927 70871
rect 36985 70825 37031 70871
rect 37089 70825 37135 70871
rect 37193 70825 37239 70871
rect 37297 70825 37343 70871
rect 37401 70825 37447 70871
rect 37505 70825 37551 70871
rect 37609 70825 37655 70871
rect 37713 70825 37759 70871
rect 37817 70825 37863 70871
rect 37921 70825 37967 70871
rect 38025 70825 38071 70871
rect 38129 70825 38175 70871
rect 38233 70825 38279 70871
rect 38337 70825 38383 70871
rect 38441 70825 38487 70871
rect 38545 70825 38591 70871
rect 38649 70825 38695 70871
rect 38753 70825 38799 70871
rect 38857 70825 38903 70871
rect 38961 70825 39007 70871
rect 39065 70825 39111 70871
rect 39169 70825 39215 70871
rect 39273 70825 39319 70871
rect 39377 70825 39423 70871
rect 39481 70825 39527 70871
rect 39585 70825 39631 70871
rect 39689 70825 39735 70871
rect 39793 70825 39839 70871
rect 39897 70825 39943 70871
rect 40001 70825 40047 70871
rect 40105 70825 40151 70871
rect 40209 70825 40255 70871
rect 40313 70825 40359 70871
rect 40417 70825 40463 70871
rect 40521 70825 40567 70871
rect 40625 70825 40671 70871
rect 40729 70825 40775 70871
rect 40833 70825 40879 70871
rect 40937 70825 40983 70871
rect 41041 70825 41087 70871
rect 41145 70825 41191 70871
rect 41249 70825 41295 70871
rect 41353 70825 41399 70871
rect 41457 70825 41503 70871
rect 41561 70825 41607 70871
rect 41665 70825 41711 70871
rect 41769 70825 41815 70871
rect 41873 70825 41919 70871
rect 41977 70825 42023 70871
rect 42081 70825 42127 70871
rect 42185 70825 42231 70871
rect 42289 70825 42335 70871
rect 42393 70825 42439 70871
rect 42497 70825 42543 70871
rect 42601 70825 42647 70871
rect 42705 70825 42751 70871
rect 42809 70825 42855 70871
rect 42913 70825 42959 70871
rect 43017 70825 43063 70871
rect 43121 70825 43167 70871
rect 43225 70825 43271 70871
rect 43329 70825 43375 70871
rect 43433 70825 43479 70871
rect 43537 70825 43583 70871
rect 43641 70825 43687 70871
rect 43745 70825 43791 70871
rect 43849 70825 43895 70871
rect 43953 70825 43999 70871
rect 44057 70825 44103 70871
rect 44161 70825 44207 70871
rect 44265 70825 44311 70871
rect 44369 70825 44415 70871
rect 44473 70825 44519 70871
rect 44577 70825 44623 70871
rect 44681 70825 44727 70871
rect 44785 70825 44831 70871
rect 44889 70825 44935 70871
rect 44993 70825 45039 70871
rect 45097 70825 45143 70871
rect 45201 70825 45247 70871
rect 45305 70825 45351 70871
rect 45409 70825 45455 70871
rect 45513 70825 45559 70871
rect 45617 70825 45663 70871
rect 45721 70825 45767 70871
rect 45825 70825 45871 70871
rect 45929 70825 45975 70871
rect 46033 70825 46079 70871
rect 46137 70825 46183 70871
rect 46241 70825 46287 70871
rect 46345 70825 46391 70871
rect 46449 70825 46495 70871
rect 46553 70825 46599 70871
rect 46657 70825 46703 70871
rect 46761 70825 46807 70871
rect 46865 70825 46911 70871
rect 46969 70825 47015 70871
rect 47073 70825 47119 70871
rect 47177 70825 47223 70871
rect 47281 70825 47327 70871
rect 47385 70825 47431 70871
rect 47489 70825 47535 70871
rect 47593 70825 47639 70871
rect 47697 70825 47743 70871
rect 47801 70825 47847 70871
rect 47905 70825 47951 70871
rect 48009 70825 48055 70871
rect 48113 70825 48159 70871
rect 48217 70825 48263 70871
rect 48321 70825 48367 70871
rect 48425 70825 48471 70871
rect 48529 70825 48575 70871
rect 48633 70825 48679 70871
rect 48737 70825 48783 70871
rect 48841 70825 48887 70871
rect 48945 70825 48991 70871
rect 49049 70825 49095 70871
rect 49153 70825 49199 70871
rect 49257 70825 49303 70871
rect 49361 70825 49407 70871
rect 49465 70825 49511 70871
rect 49569 70825 49615 70871
rect 49673 70825 49719 70871
rect 49777 70825 49823 70871
rect 49881 70825 49927 70871
rect 49985 70825 50031 70871
rect 50089 70825 50135 70871
rect 50193 70825 50239 70871
rect 50297 70825 50343 70871
rect 50401 70825 50447 70871
rect 50505 70825 50551 70871
rect 50609 70825 50655 70871
rect 50713 70825 50759 70871
rect 50817 70825 50863 70871
rect 50921 70825 50967 70871
rect 51025 70825 51071 70871
rect 51129 70825 51175 70871
rect 51233 70825 51279 70871
rect 51337 70825 51383 70871
rect 51441 70825 51487 70871
rect 51545 70825 51591 70871
rect 51649 70825 51695 70871
rect 51753 70825 51799 70871
rect 51857 70825 51903 70871
rect 51961 70825 52007 70871
rect 52065 70825 52111 70871
rect 52169 70825 52215 70871
rect 52273 70825 52319 70871
rect 52377 70825 52423 70871
rect 52481 70825 52527 70871
rect 52585 70825 52631 70871
rect 52689 70825 52735 70871
rect 52793 70825 52839 70871
rect 52897 70825 52943 70871
rect 53001 70825 53047 70871
rect 53105 70825 53151 70871
rect 53209 70825 53255 70871
rect 53313 70825 53359 70871
rect 53417 70825 53463 70871
rect 53521 70825 53567 70871
rect 53625 70825 53671 70871
rect 53729 70825 53775 70871
rect 53833 70825 53879 70871
rect 53937 70825 53983 70871
rect 54041 70825 54087 70871
rect 54145 70825 54191 70871
rect 54249 70825 54295 70871
rect 54353 70825 54399 70871
rect 54457 70825 54503 70871
rect 54561 70825 54607 70871
rect 54665 70825 54711 70871
rect 54769 70825 54815 70871
rect 54873 70825 54919 70871
rect 54977 70825 55023 70871
rect 55081 70825 55127 70871
rect 55185 70825 55231 70871
rect 55289 70825 55335 70871
rect 55393 70825 55439 70871
rect 55497 70825 55543 70871
rect 55601 70825 55647 70871
rect 55705 70825 55751 70871
rect 55809 70825 55855 70871
rect 55913 70825 55959 70871
rect 56017 70825 56063 70871
rect 56121 70825 56167 70871
rect 56225 70825 56271 70871
rect 56329 70825 56375 70871
rect 56433 70825 56479 70871
rect 56537 70825 56583 70871
rect 56641 70825 56687 70871
rect 56745 70825 56791 70871
rect 56849 70825 56895 70871
rect 56953 70825 56999 70871
rect 57057 70825 57103 70871
rect 57161 70825 57207 70871
rect 57265 70825 57311 70871
rect 57369 70825 57415 70871
rect 57473 70825 57519 70871
rect 57577 70825 57623 70871
rect 57681 70825 57727 70871
rect 57785 70825 57831 70871
rect 57889 70825 57935 70871
rect 57993 70825 58039 70871
rect 58097 70825 58143 70871
rect 58201 70825 58247 70871
rect 58305 70825 58351 70871
rect 58409 70825 58455 70871
rect 58513 70825 58559 70871
rect 58617 70825 58663 70871
rect 58721 70825 58767 70871
rect 58825 70825 58871 70871
rect 58929 70825 58975 70871
rect 59033 70825 59079 70871
rect 59137 70825 59183 70871
rect 59241 70825 59287 70871
rect 59345 70825 59391 70871
rect 59449 70825 59495 70871
rect 59553 70825 59599 70871
rect 59657 70825 59703 70871
rect 59761 70825 59807 70871
rect 59865 70825 59911 70871
rect 59969 70825 60015 70871
rect 60073 70825 60119 70871
rect 60177 70825 60223 70871
rect 60281 70825 60327 70871
rect 60385 70825 60431 70871
rect 60489 70825 60535 70871
rect 60593 70825 60639 70871
rect 60697 70825 60743 70871
rect 60801 70825 60847 70871
rect 60905 70825 60951 70871
rect 61009 70825 61055 70871
rect 61113 70825 61159 70871
rect 61217 70825 61263 70871
rect 61321 70825 61367 70871
rect 61425 70825 61471 70871
rect 61529 70825 61575 70871
rect 61633 70825 61679 70871
rect 61737 70825 61783 70871
rect 61841 70825 61887 70871
rect 61945 70825 61991 70871
rect 62049 70825 62095 70871
rect 62153 70825 62199 70871
rect 62257 70825 62303 70871
rect 62361 70825 62407 70871
rect 62465 70825 62511 70871
rect 62569 70825 62615 70871
rect 62673 70825 62719 70871
rect 62777 70825 62823 70871
rect 62881 70825 62927 70871
rect 62985 70825 63031 70871
rect 63089 70825 63135 70871
rect 63193 70825 63239 70871
rect 63297 70825 63343 70871
rect 63401 70825 63447 70871
rect 63505 70825 63551 70871
rect 63609 70825 63655 70871
rect 63713 70825 63759 70871
rect 63817 70825 63863 70871
rect 63921 70825 63967 70871
rect 64025 70825 64071 70871
rect 64129 70825 64175 70871
rect 64233 70825 64279 70871
rect 64337 70825 64383 70871
rect 64441 70825 64487 70871
rect 64545 70825 64591 70871
rect 64649 70825 64695 70871
rect 64753 70825 64799 70871
rect 64857 70825 64903 70871
rect 64961 70825 65007 70871
rect 65065 70825 65111 70871
rect 65169 70825 65215 70871
rect 65273 70825 65319 70871
rect 65377 70825 65423 70871
rect 65481 70825 65527 70871
rect 65585 70825 65631 70871
rect 65689 70825 65735 70871
rect 65793 70825 65839 70871
rect 65897 70825 65943 70871
rect 66001 70825 66047 70871
rect 66105 70825 66151 70871
rect 66209 70825 66255 70871
rect 66313 70825 66359 70871
rect 66417 70825 66463 70871
rect 66521 70825 66567 70871
rect 66625 70825 66671 70871
rect 66729 70825 66775 70871
rect 66833 70825 66879 70871
rect 66937 70825 66983 70871
rect 67041 70825 67087 70871
rect 67145 70825 67191 70871
rect 67249 70825 67295 70871
rect 67353 70825 67399 70871
rect 67457 70825 67503 70871
rect 67561 70825 67607 70871
rect 67665 70825 67711 70871
rect 67769 70825 67815 70871
rect 67873 70825 67919 70871
rect 67977 70825 68023 70871
rect 68081 70825 68127 70871
rect 68185 70825 68231 70871
rect 68289 70825 68335 70871
rect 68393 70825 68439 70871
rect 68497 70825 68543 70871
rect 68601 70825 68647 70871
rect 68705 70825 68751 70871
rect 68809 70825 68855 70871
rect 68913 70825 68959 70871
rect 69017 70825 69063 70871
rect 69121 70825 69167 70871
rect 69225 70825 69271 70871
rect 69329 70825 69375 70871
rect 69433 70825 69479 70871
rect 69537 70825 69583 70871
rect 69641 70825 69687 70871
rect 69745 70825 69791 70871
rect 69849 70825 69895 70871
rect 13119 70721 13165 70767
rect 13223 70721 13269 70767
rect 13119 70617 13165 70663
rect 13223 70617 13269 70663
rect 13119 70513 13165 70559
rect 13223 70513 13269 70559
rect 13119 70409 13165 70455
rect 13223 70409 13269 70455
rect 13119 70305 13165 70351
rect 13223 70305 13269 70351
rect 13119 70201 13165 70247
rect 13223 70201 13269 70247
rect 13119 70097 13165 70143
rect 13223 70097 13269 70143
rect 13119 69993 13165 70039
rect 13223 69993 13269 70039
rect 13119 69889 13165 69935
rect 13223 69889 13269 69935
rect 13119 69785 13165 69831
rect 13223 69785 13269 69831
rect 69796 70674 69842 70720
rect 69900 70674 69946 70720
rect 69796 70570 69842 70616
rect 69900 70570 69946 70616
rect 69796 70466 69842 70512
rect 69900 70466 69946 70512
rect 69796 70362 69842 70408
rect 69900 70362 69946 70408
rect 69796 70258 69842 70304
rect 69900 70258 69946 70304
rect 69796 70154 69842 70200
rect 69900 70154 69946 70200
rect 69796 70050 69842 70096
rect 69900 70050 69946 70096
rect 69796 69900 69842 69946
rect 69900 69900 69946 69946
rect 70004 69900 70050 69946
rect 70108 69900 70154 69946
rect 70212 69900 70258 69946
rect 70316 69900 70362 69946
rect 70420 69900 70466 69946
rect 70524 69900 70570 69946
rect 70628 69900 70674 69946
rect 70824 69862 70870 69908
rect 70928 69862 70974 69908
rect 69796 69796 69842 69842
rect 69900 69796 69946 69842
rect 70004 69796 70050 69842
rect 70108 69796 70154 69842
rect 70212 69796 70258 69842
rect 70316 69796 70362 69842
rect 70420 69796 70466 69842
rect 70524 69796 70570 69842
rect 70628 69796 70674 69842
rect 13119 69681 13165 69727
rect 13223 69681 13269 69727
rect 13119 69577 13165 69623
rect 13223 69577 13269 69623
rect 13119 69473 13165 69519
rect 13223 69473 13269 69519
rect 13119 69369 13165 69415
rect 13223 69369 13269 69415
rect 13119 69265 13165 69311
rect 13223 69265 13269 69311
rect 13119 69161 13165 69207
rect 13223 69161 13269 69207
rect 13119 69057 13165 69103
rect 13223 69057 13269 69103
rect 13119 68953 13165 68999
rect 13223 68953 13269 68999
rect 13119 68849 13165 68895
rect 13223 68849 13269 68895
rect 13119 68745 13165 68791
rect 13223 68745 13269 68791
rect 13119 68641 13165 68687
rect 13223 68641 13269 68687
rect 13119 68537 13165 68583
rect 13223 68537 13269 68583
rect 13119 68433 13165 68479
rect 13223 68433 13269 68479
rect 13119 68329 13165 68375
rect 13223 68329 13269 68375
rect 13119 68225 13165 68271
rect 13223 68225 13269 68271
rect 13119 68121 13165 68167
rect 13223 68121 13269 68167
rect 13119 68017 13165 68063
rect 13223 68017 13269 68063
rect 13119 67913 13165 67959
rect 13223 67913 13269 67959
rect 13119 67809 13165 67855
rect 13223 67809 13269 67855
rect 13119 67705 13165 67751
rect 13223 67705 13269 67751
rect 13119 67601 13165 67647
rect 13223 67601 13269 67647
rect 13119 67497 13165 67543
rect 13223 67497 13269 67543
rect 13119 67393 13165 67439
rect 13223 67393 13269 67439
rect 13119 67289 13165 67335
rect 13223 67289 13269 67335
rect 13119 67185 13165 67231
rect 13223 67185 13269 67231
rect 13119 67081 13165 67127
rect 13223 67081 13269 67127
rect 13119 66977 13165 67023
rect 13223 66977 13269 67023
rect 13119 66873 13165 66919
rect 13223 66873 13269 66919
rect 13119 66769 13165 66815
rect 13223 66769 13269 66815
rect 13119 66665 13165 66711
rect 13223 66665 13269 66711
rect 13119 66561 13165 66607
rect 13223 66561 13269 66607
rect 13119 66457 13165 66503
rect 13223 66457 13269 66503
rect 13119 66353 13165 66399
rect 13223 66353 13269 66399
rect 13119 66249 13165 66295
rect 13223 66249 13269 66295
rect 13119 66145 13165 66191
rect 13223 66145 13269 66191
rect 13119 66041 13165 66087
rect 13223 66041 13269 66087
rect 13119 65937 13165 65983
rect 13223 65937 13269 65983
rect 13119 65833 13165 65879
rect 13223 65833 13269 65879
rect 13119 65729 13165 65775
rect 13223 65729 13269 65775
rect 13119 65625 13165 65671
rect 13223 65625 13269 65671
rect 13119 65521 13165 65567
rect 13223 65521 13269 65567
rect 13119 65417 13165 65463
rect 13223 65417 13269 65463
rect 13119 65313 13165 65359
rect 13223 65313 13269 65359
rect 13119 65209 13165 65255
rect 13223 65209 13269 65255
rect 13119 65105 13165 65151
rect 13223 65105 13269 65151
rect 13119 65001 13165 65047
rect 13223 65001 13269 65047
rect 13119 64897 13165 64943
rect 13223 64897 13269 64943
rect 13119 64793 13165 64839
rect 13223 64793 13269 64839
rect 13119 64689 13165 64735
rect 13223 64689 13269 64735
rect 13119 64585 13165 64631
rect 13223 64585 13269 64631
rect 13119 64481 13165 64527
rect 13223 64481 13269 64527
rect 13119 64377 13165 64423
rect 13223 64377 13269 64423
rect 13119 64273 13165 64319
rect 13223 64273 13269 64319
rect 13119 64169 13165 64215
rect 13223 64169 13269 64215
rect 13119 64065 13165 64111
rect 13223 64065 13269 64111
rect 13119 63961 13165 64007
rect 13223 63961 13269 64007
rect 13119 63857 13165 63903
rect 13223 63857 13269 63903
rect 13119 63753 13165 63799
rect 13223 63753 13269 63799
rect 13119 63649 13165 63695
rect 13223 63649 13269 63695
rect 13119 63545 13165 63591
rect 13223 63545 13269 63591
rect 13119 63441 13165 63487
rect 13223 63441 13269 63487
rect 13119 63337 13165 63383
rect 13223 63337 13269 63383
rect 13119 63233 13165 63279
rect 13223 63233 13269 63279
rect 13119 63129 13165 63175
rect 13223 63129 13269 63175
rect 13119 63025 13165 63071
rect 13223 63025 13269 63071
rect 13119 62921 13165 62967
rect 13223 62921 13269 62967
rect 13119 62817 13165 62863
rect 13223 62817 13269 62863
rect 13119 62713 13165 62759
rect 13223 62713 13269 62759
rect 13119 62609 13165 62655
rect 13223 62609 13269 62655
rect 13119 62505 13165 62551
rect 13223 62505 13269 62551
rect 13119 62401 13165 62447
rect 13223 62401 13269 62447
rect 13119 62297 13165 62343
rect 13223 62297 13269 62343
rect 13119 62193 13165 62239
rect 13223 62193 13269 62239
rect 13119 62089 13165 62135
rect 13223 62089 13269 62135
rect 13119 61985 13165 62031
rect 13223 61985 13269 62031
rect 13119 61881 13165 61927
rect 13223 61881 13269 61927
rect 13119 61777 13165 61823
rect 13223 61777 13269 61823
rect 13119 61673 13165 61719
rect 13223 61673 13269 61719
rect 13119 61569 13165 61615
rect 13223 61569 13269 61615
rect 13119 61465 13165 61511
rect 13223 61465 13269 61511
rect 13119 61361 13165 61407
rect 13223 61361 13269 61407
rect 13119 61257 13165 61303
rect 13223 61257 13269 61303
rect 13119 61153 13165 61199
rect 13223 61153 13269 61199
rect 13119 61049 13165 61095
rect 13223 61049 13269 61095
rect 13119 60945 13165 60991
rect 13223 60945 13269 60991
rect 13119 60841 13165 60887
rect 13223 60841 13269 60887
rect 13119 60737 13165 60783
rect 13223 60737 13269 60783
rect 13119 60633 13165 60679
rect 13223 60633 13269 60679
rect 13119 60529 13165 60575
rect 13223 60529 13269 60575
rect 13119 60425 13165 60471
rect 13223 60425 13269 60471
rect 13119 60321 13165 60367
rect 13223 60321 13269 60367
rect 13119 60217 13165 60263
rect 13223 60217 13269 60263
rect 13119 60113 13165 60159
rect 13223 60113 13269 60159
rect 13119 60009 13165 60055
rect 13223 60009 13269 60055
rect 13119 59905 13165 59951
rect 13223 59905 13269 59951
rect 13119 59801 13165 59847
rect 13223 59801 13269 59847
rect 13119 59697 13165 59743
rect 13223 59697 13269 59743
rect 13119 59593 13165 59639
rect 13223 59593 13269 59639
rect 13119 59489 13165 59535
rect 13223 59489 13269 59535
rect 13119 59385 13165 59431
rect 13223 59385 13269 59431
rect 13119 59281 13165 59327
rect 13223 59281 13269 59327
rect 13119 59177 13165 59223
rect 13223 59177 13269 59223
rect 13119 59073 13165 59119
rect 13223 59073 13269 59119
rect 13119 58969 13165 59015
rect 13223 58969 13269 59015
rect 13119 58865 13165 58911
rect 13223 58865 13269 58911
rect 13119 58761 13165 58807
rect 13223 58761 13269 58807
rect 13119 58657 13165 58703
rect 13223 58657 13269 58703
rect 13119 58553 13165 58599
rect 13223 58553 13269 58599
rect 13119 58449 13165 58495
rect 13223 58449 13269 58495
rect 13119 58345 13165 58391
rect 13223 58345 13269 58391
rect 13119 58241 13165 58287
rect 13223 58241 13269 58287
rect 13119 58137 13165 58183
rect 13223 58137 13269 58183
rect 13119 58033 13165 58079
rect 13223 58033 13269 58079
rect 13119 57929 13165 57975
rect 13223 57929 13269 57975
rect 13119 57825 13165 57871
rect 13223 57825 13269 57871
rect 13119 57721 13165 57767
rect 13223 57721 13269 57767
rect 13119 57617 13165 57663
rect 13223 57617 13269 57663
rect 13119 57513 13165 57559
rect 13223 57513 13269 57559
rect 13119 57409 13165 57455
rect 13223 57409 13269 57455
rect 13119 57305 13165 57351
rect 13223 57305 13269 57351
rect 13119 57201 13165 57247
rect 13223 57201 13269 57247
rect 13119 57097 13165 57143
rect 13223 57097 13269 57143
rect 13119 56993 13165 57039
rect 13223 56993 13269 57039
rect 13119 56889 13165 56935
rect 13223 56889 13269 56935
rect 13119 56785 13165 56831
rect 13223 56785 13269 56831
rect 13119 56681 13165 56727
rect 13223 56681 13269 56727
rect 13119 56577 13165 56623
rect 13223 56577 13269 56623
rect 13119 56473 13165 56519
rect 13223 56473 13269 56519
rect 13119 56369 13165 56415
rect 13223 56369 13269 56415
rect 13119 56265 13165 56311
rect 13223 56265 13269 56311
rect 13119 56161 13165 56207
rect 13223 56161 13269 56207
rect 13119 56057 13165 56103
rect 13223 56057 13269 56103
rect 13119 55953 13165 55999
rect 13223 55953 13269 55999
rect 13119 55849 13165 55895
rect 13223 55849 13269 55895
rect 13119 55745 13165 55791
rect 13223 55745 13269 55791
rect 13119 55641 13165 55687
rect 13223 55641 13269 55687
rect 13119 55537 13165 55583
rect 13223 55537 13269 55583
rect 13119 55433 13165 55479
rect 13223 55433 13269 55479
rect 13119 55329 13165 55375
rect 13223 55329 13269 55375
rect 13119 55225 13165 55271
rect 13223 55225 13269 55271
rect 13119 55121 13165 55167
rect 13223 55121 13269 55167
rect 13119 55017 13165 55063
rect 13223 55017 13269 55063
rect 13119 54913 13165 54959
rect 13223 54913 13269 54959
rect 13119 54809 13165 54855
rect 13223 54809 13269 54855
rect 13119 54705 13165 54751
rect 13223 54705 13269 54751
rect 13119 54601 13165 54647
rect 13223 54601 13269 54647
rect 13119 54497 13165 54543
rect 13223 54497 13269 54543
rect 13119 54393 13165 54439
rect 13223 54393 13269 54439
rect 13119 54289 13165 54335
rect 13223 54289 13269 54335
rect 13119 54185 13165 54231
rect 13223 54185 13269 54231
rect 13119 54081 13165 54127
rect 13223 54081 13269 54127
rect 13119 53977 13165 54023
rect 13223 53977 13269 54023
rect 13119 53873 13165 53919
rect 13223 53873 13269 53919
rect 13119 53769 13165 53815
rect 13223 53769 13269 53815
rect 13119 53665 13165 53711
rect 13223 53665 13269 53711
rect 13119 53561 13165 53607
rect 13223 53561 13269 53607
rect 13119 53457 13165 53503
rect 13223 53457 13269 53503
rect 13119 53353 13165 53399
rect 13223 53353 13269 53399
rect 13119 53249 13165 53295
rect 13223 53249 13269 53295
rect 13119 53145 13165 53191
rect 13223 53145 13269 53191
rect 13119 53041 13165 53087
rect 13223 53041 13269 53087
rect 13119 52937 13165 52983
rect 13223 52937 13269 52983
rect 13119 52833 13165 52879
rect 13223 52833 13269 52879
rect 13119 52729 13165 52775
rect 13223 52729 13269 52775
rect 13119 52625 13165 52671
rect 13223 52625 13269 52671
rect 13119 52521 13165 52567
rect 13223 52521 13269 52567
rect 13119 52417 13165 52463
rect 13223 52417 13269 52463
rect 13119 52313 13165 52359
rect 13223 52313 13269 52359
rect 13119 52209 13165 52255
rect 13223 52209 13269 52255
rect 13119 52105 13165 52151
rect 13223 52105 13269 52151
rect 13119 52001 13165 52047
rect 13223 52001 13269 52047
rect 13119 51897 13165 51943
rect 13223 51897 13269 51943
rect 13119 51793 13165 51839
rect 13223 51793 13269 51839
rect 13119 51689 13165 51735
rect 13223 51689 13269 51735
rect 13119 51585 13165 51631
rect 13223 51585 13269 51631
rect 13119 51481 13165 51527
rect 13223 51481 13269 51527
rect 13119 51377 13165 51423
rect 13223 51377 13269 51423
rect 13119 51273 13165 51319
rect 13223 51273 13269 51319
rect 13119 51169 13165 51215
rect 13223 51169 13269 51215
rect 13119 51065 13165 51111
rect 13223 51065 13269 51111
rect 13119 50961 13165 51007
rect 13223 50961 13269 51007
rect 13119 50857 13165 50903
rect 13223 50857 13269 50903
rect 13119 50753 13165 50799
rect 13223 50753 13269 50799
rect 13119 50649 13165 50695
rect 13223 50649 13269 50695
rect 13119 50545 13165 50591
rect 13223 50545 13269 50591
rect 13119 50441 13165 50487
rect 13223 50441 13269 50487
rect 13119 50337 13165 50383
rect 13223 50337 13269 50383
rect 13119 50233 13165 50279
rect 13223 50233 13269 50279
rect 13119 50129 13165 50175
rect 13223 50129 13269 50175
rect 13119 50025 13165 50071
rect 13223 50025 13269 50071
rect 13119 49921 13165 49967
rect 13223 49921 13269 49967
rect 13119 49817 13165 49863
rect 13223 49817 13269 49863
rect 13119 49713 13165 49759
rect 13223 49713 13269 49759
rect 13119 49609 13165 49655
rect 13223 49609 13269 49655
rect 13119 49505 13165 49551
rect 13223 49505 13269 49551
rect 13119 49401 13165 49447
rect 13223 49401 13269 49447
rect 13119 49297 13165 49343
rect 13223 49297 13269 49343
rect 13119 49193 13165 49239
rect 13223 49193 13269 49239
rect 13119 49089 13165 49135
rect 13223 49089 13269 49135
rect 13119 48985 13165 49031
rect 13223 48985 13269 49031
rect 13119 48881 13165 48927
rect 13223 48881 13269 48927
rect 13119 48777 13165 48823
rect 13223 48777 13269 48823
rect 13119 48673 13165 48719
rect 13223 48673 13269 48719
rect 13119 48569 13165 48615
rect 13223 48569 13269 48615
rect 13119 48465 13165 48511
rect 13223 48465 13269 48511
rect 13119 48361 13165 48407
rect 13223 48361 13269 48407
rect 13119 48257 13165 48303
rect 13223 48257 13269 48303
rect 13119 48153 13165 48199
rect 13223 48153 13269 48199
rect 13119 48049 13165 48095
rect 13223 48049 13269 48095
rect 13119 47945 13165 47991
rect 13223 47945 13269 47991
rect 13119 47841 13165 47887
rect 13223 47841 13269 47887
rect 13119 47737 13165 47783
rect 13223 47737 13269 47783
rect 13119 47633 13165 47679
rect 13223 47633 13269 47679
rect 13119 47529 13165 47575
rect 13223 47529 13269 47575
rect 13119 47425 13165 47471
rect 13223 47425 13269 47471
rect 13119 47321 13165 47367
rect 13223 47321 13269 47367
rect 13119 47217 13165 47263
rect 13223 47217 13269 47263
rect 13119 47113 13165 47159
rect 13223 47113 13269 47159
rect 13119 47009 13165 47055
rect 13223 47009 13269 47055
rect 13119 46905 13165 46951
rect 13223 46905 13269 46951
rect 13119 46801 13165 46847
rect 13223 46801 13269 46847
rect 13119 46697 13165 46743
rect 13223 46697 13269 46743
rect 13119 46593 13165 46639
rect 13223 46593 13269 46639
rect 13119 46489 13165 46535
rect 13223 46489 13269 46535
rect 13119 46385 13165 46431
rect 13223 46385 13269 46431
rect 13119 46281 13165 46327
rect 13223 46281 13269 46327
rect 13119 46177 13165 46223
rect 13223 46177 13269 46223
rect 13119 46073 13165 46119
rect 13223 46073 13269 46119
rect 13119 45969 13165 46015
rect 13223 45969 13269 46015
rect 13119 45865 13165 45911
rect 13223 45865 13269 45911
rect 13119 45761 13165 45807
rect 13223 45761 13269 45807
rect 13119 45657 13165 45703
rect 13223 45657 13269 45703
rect 13119 45553 13165 45599
rect 13223 45553 13269 45599
rect 13119 45449 13165 45495
rect 13223 45449 13269 45495
rect 13119 45345 13165 45391
rect 13223 45345 13269 45391
rect 13119 45241 13165 45287
rect 13223 45241 13269 45287
rect 13119 45137 13165 45183
rect 13223 45137 13269 45183
rect 13119 45033 13165 45079
rect 13223 45033 13269 45079
rect 70824 69758 70870 69804
rect 70928 69758 70974 69804
rect 70824 69654 70870 69700
rect 70928 69654 70974 69700
rect 70824 69550 70870 69596
rect 70928 69550 70974 69596
rect 70824 69446 70870 69492
rect 70928 69446 70974 69492
rect 70824 69342 70870 69388
rect 70928 69342 70974 69388
rect 70824 69238 70870 69284
rect 70928 69238 70974 69284
rect 70824 69134 70870 69180
rect 70928 69134 70974 69180
rect 70824 69030 70870 69076
rect 70928 69030 70974 69076
rect 70824 68926 70870 68972
rect 70928 68926 70974 68972
rect 70824 68822 70870 68868
rect 70928 68822 70974 68868
rect 70824 68718 70870 68764
rect 70928 68718 70974 68764
rect 70824 68614 70870 68660
rect 70928 68614 70974 68660
rect 70824 68510 70870 68556
rect 70928 68510 70974 68556
rect 70824 68406 70870 68452
rect 70928 68406 70974 68452
rect 70824 68302 70870 68348
rect 70928 68302 70974 68348
rect 70824 68198 70870 68244
rect 70928 68198 70974 68244
rect 70824 68094 70870 68140
rect 70928 68094 70974 68140
rect 70824 67990 70870 68036
rect 70928 67990 70974 68036
rect 70824 67886 70870 67932
rect 70928 67886 70974 67932
rect 70824 67782 70870 67828
rect 70928 67782 70974 67828
rect 70824 67678 70870 67724
rect 70928 67678 70974 67724
rect 70824 67574 70870 67620
rect 70928 67574 70974 67620
rect 70824 67470 70870 67516
rect 70928 67470 70974 67516
rect 70824 67366 70870 67412
rect 70928 67366 70974 67412
rect 70824 67262 70870 67308
rect 70928 67262 70974 67308
rect 70824 67158 70870 67204
rect 70928 67158 70974 67204
rect 70824 67054 70870 67100
rect 70928 67054 70974 67100
rect 70824 66950 70870 66996
rect 70928 66950 70974 66996
rect 70824 66846 70870 66892
rect 70928 66846 70974 66892
rect 70824 66742 70870 66788
rect 70928 66742 70974 66788
rect 70824 66638 70870 66684
rect 70928 66638 70974 66684
rect 70824 66534 70870 66580
rect 70928 66534 70974 66580
rect 70824 66430 70870 66476
rect 70928 66430 70974 66476
rect 70824 66326 70870 66372
rect 70928 66326 70974 66372
rect 70824 66222 70870 66268
rect 70928 66222 70974 66268
rect 70824 66118 70870 66164
rect 70928 66118 70974 66164
rect 70824 66014 70870 66060
rect 70928 66014 70974 66060
rect 70824 65910 70870 65956
rect 70928 65910 70974 65956
rect 70824 65806 70870 65852
rect 70928 65806 70974 65852
rect 70824 65702 70870 65748
rect 70928 65702 70974 65748
rect 70824 65598 70870 65644
rect 70928 65598 70974 65644
rect 70824 65494 70870 65540
rect 70928 65494 70974 65540
rect 70824 65390 70870 65436
rect 70928 65390 70974 65436
rect 70824 65286 70870 65332
rect 70928 65286 70974 65332
rect 70824 65182 70870 65228
rect 70928 65182 70974 65228
rect 70824 65078 70870 65124
rect 70928 65078 70974 65124
rect 70824 64974 70870 65020
rect 70928 64974 70974 65020
rect 70824 64870 70870 64916
rect 70928 64870 70974 64916
rect 70824 64766 70870 64812
rect 70928 64766 70974 64812
rect 70824 64662 70870 64708
rect 70928 64662 70974 64708
rect 70824 64558 70870 64604
rect 70928 64558 70974 64604
rect 70824 64454 70870 64500
rect 70928 64454 70974 64500
rect 70824 64350 70870 64396
rect 70928 64350 70974 64396
rect 70824 64246 70870 64292
rect 70928 64246 70974 64292
rect 70824 64142 70870 64188
rect 70928 64142 70974 64188
rect 70824 64038 70870 64084
rect 70928 64038 70974 64084
rect 70824 63934 70870 63980
rect 70928 63934 70974 63980
rect 70824 63830 70870 63876
rect 70928 63830 70974 63876
rect 70824 63726 70870 63772
rect 70928 63726 70974 63772
rect 70824 63622 70870 63668
rect 70928 63622 70974 63668
rect 70824 63518 70870 63564
rect 70928 63518 70974 63564
rect 70824 63414 70870 63460
rect 70928 63414 70974 63460
rect 70824 63310 70870 63356
rect 70928 63310 70974 63356
rect 70824 63206 70870 63252
rect 70928 63206 70974 63252
rect 70824 63102 70870 63148
rect 70928 63102 70974 63148
rect 70824 62998 70870 63044
rect 70928 62998 70974 63044
rect 70824 62894 70870 62940
rect 70928 62894 70974 62940
rect 70824 62790 70870 62836
rect 70928 62790 70974 62836
rect 70824 62686 70870 62732
rect 70928 62686 70974 62732
rect 70824 62582 70870 62628
rect 70928 62582 70974 62628
rect 70824 62478 70870 62524
rect 70928 62478 70974 62524
rect 70824 62374 70870 62420
rect 70928 62374 70974 62420
rect 70824 62270 70870 62316
rect 70928 62270 70974 62316
rect 70824 62166 70870 62212
rect 70928 62166 70974 62212
rect 70824 62062 70870 62108
rect 70928 62062 70974 62108
rect 70824 61958 70870 62004
rect 70928 61958 70974 62004
rect 70824 61854 70870 61900
rect 70928 61854 70974 61900
rect 70824 61750 70870 61796
rect 70928 61750 70974 61796
rect 70824 61646 70870 61692
rect 70928 61646 70974 61692
rect 70824 61542 70870 61588
rect 70928 61542 70974 61588
rect 70824 61438 70870 61484
rect 70928 61438 70974 61484
rect 70824 61334 70870 61380
rect 70928 61334 70974 61380
rect 70824 61230 70870 61276
rect 70928 61230 70974 61276
rect 70824 61126 70870 61172
rect 70928 61126 70974 61172
rect 70824 61022 70870 61068
rect 70928 61022 70974 61068
rect 70824 60918 70870 60964
rect 70928 60918 70974 60964
rect 70824 60814 70870 60860
rect 70928 60814 70974 60860
rect 70824 60710 70870 60756
rect 70928 60710 70974 60756
rect 70824 60606 70870 60652
rect 70928 60606 70974 60652
rect 70824 60502 70870 60548
rect 70928 60502 70974 60548
rect 70824 60398 70870 60444
rect 70928 60398 70974 60444
rect 70824 60294 70870 60340
rect 70928 60294 70974 60340
rect 70824 60190 70870 60236
rect 70928 60190 70974 60236
rect 70824 60086 70870 60132
rect 70928 60086 70974 60132
rect 70824 59982 70870 60028
rect 70928 59982 70974 60028
rect 70824 59878 70870 59924
rect 70928 59878 70974 59924
rect 70824 59774 70870 59820
rect 70928 59774 70974 59820
rect 70824 59670 70870 59716
rect 70928 59670 70974 59716
rect 70824 59566 70870 59612
rect 70928 59566 70974 59612
rect 70824 59462 70870 59508
rect 70928 59462 70974 59508
rect 70824 59358 70870 59404
rect 70928 59358 70974 59404
rect 70824 59254 70870 59300
rect 70928 59254 70974 59300
rect 70824 59150 70870 59196
rect 70928 59150 70974 59196
rect 70824 59046 70870 59092
rect 70928 59046 70974 59092
rect 70824 58942 70870 58988
rect 70928 58942 70974 58988
rect 70824 58838 70870 58884
rect 70928 58838 70974 58884
rect 70824 58734 70870 58780
rect 70928 58734 70974 58780
rect 70824 58630 70870 58676
rect 70928 58630 70974 58676
rect 70824 58526 70870 58572
rect 70928 58526 70974 58572
rect 70824 58422 70870 58468
rect 70928 58422 70974 58468
rect 70824 58318 70870 58364
rect 70928 58318 70974 58364
rect 70824 58214 70870 58260
rect 70928 58214 70974 58260
rect 70824 58110 70870 58156
rect 70928 58110 70974 58156
rect 70824 58006 70870 58052
rect 70928 58006 70974 58052
rect 70824 57902 70870 57948
rect 70928 57902 70974 57948
rect 70824 57798 70870 57844
rect 70928 57798 70974 57844
rect 70824 57694 70870 57740
rect 70928 57694 70974 57740
rect 70824 57590 70870 57636
rect 70928 57590 70974 57636
rect 70824 57486 70870 57532
rect 70928 57486 70974 57532
rect 70824 57382 70870 57428
rect 70928 57382 70974 57428
rect 70824 57278 70870 57324
rect 70928 57278 70974 57324
rect 70824 57174 70870 57220
rect 70928 57174 70974 57220
rect 70824 57070 70870 57116
rect 70928 57070 70974 57116
rect 70824 56966 70870 57012
rect 70928 56966 70974 57012
rect 70824 56862 70870 56908
rect 70928 56862 70974 56908
rect 70824 56758 70870 56804
rect 70928 56758 70974 56804
rect 70824 56654 70870 56700
rect 70928 56654 70974 56700
rect 70824 56550 70870 56596
rect 70928 56550 70974 56596
rect 70824 56446 70870 56492
rect 70928 56446 70974 56492
rect 70824 56342 70870 56388
rect 70928 56342 70974 56388
rect 70824 56238 70870 56284
rect 70928 56238 70974 56284
rect 70824 56134 70870 56180
rect 70928 56134 70974 56180
rect 70824 56030 70870 56076
rect 70928 56030 70974 56076
rect 70824 55926 70870 55972
rect 70928 55926 70974 55972
rect 70824 55822 70870 55868
rect 70928 55822 70974 55868
rect 70824 55718 70870 55764
rect 70928 55718 70974 55764
rect 70824 55614 70870 55660
rect 70928 55614 70974 55660
rect 70824 55510 70870 55556
rect 70928 55510 70974 55556
rect 70824 55406 70870 55452
rect 70928 55406 70974 55452
rect 70824 55302 70870 55348
rect 70928 55302 70974 55348
rect 70824 55198 70870 55244
rect 70928 55198 70974 55244
rect 70824 55094 70870 55140
rect 70928 55094 70974 55140
rect 70824 54990 70870 55036
rect 70928 54990 70974 55036
rect 70824 54886 70870 54932
rect 70928 54886 70974 54932
rect 70824 54782 70870 54828
rect 70928 54782 70974 54828
rect 70824 54678 70870 54724
rect 70928 54678 70974 54724
rect 70824 54574 70870 54620
rect 70928 54574 70974 54620
rect 70824 54470 70870 54516
rect 70928 54470 70974 54516
rect 70824 54366 70870 54412
rect 70928 54366 70974 54412
rect 70824 54262 70870 54308
rect 70928 54262 70974 54308
rect 70824 54158 70870 54204
rect 70928 54158 70974 54204
rect 70824 54054 70870 54100
rect 70928 54054 70974 54100
rect 70824 53950 70870 53996
rect 70928 53950 70974 53996
rect 70824 53846 70870 53892
rect 70928 53846 70974 53892
rect 70824 53742 70870 53788
rect 70928 53742 70974 53788
rect 70824 53638 70870 53684
rect 70928 53638 70974 53684
rect 70824 53534 70870 53580
rect 70928 53534 70974 53580
rect 70824 53430 70870 53476
rect 70928 53430 70974 53476
rect 70824 53326 70870 53372
rect 70928 53326 70974 53372
rect 70824 53222 70870 53268
rect 70928 53222 70974 53268
rect 70824 53118 70870 53164
rect 70928 53118 70974 53164
rect 70824 53014 70870 53060
rect 70928 53014 70974 53060
rect 70824 52910 70870 52956
rect 70928 52910 70974 52956
rect 70824 52806 70870 52852
rect 70928 52806 70974 52852
rect 70824 52702 70870 52748
rect 70928 52702 70974 52748
rect 70824 52598 70870 52644
rect 70928 52598 70974 52644
rect 70824 52494 70870 52540
rect 70928 52494 70974 52540
rect 70824 52390 70870 52436
rect 70928 52390 70974 52436
rect 70824 52286 70870 52332
rect 70928 52286 70974 52332
rect 70824 52182 70870 52228
rect 70928 52182 70974 52228
rect 70824 52078 70870 52124
rect 70928 52078 70974 52124
rect 70824 51974 70870 52020
rect 70928 51974 70974 52020
rect 70824 51870 70870 51916
rect 70928 51870 70974 51916
rect 70824 51766 70870 51812
rect 70928 51766 70974 51812
rect 70824 51662 70870 51708
rect 70928 51662 70974 51708
rect 70824 51558 70870 51604
rect 70928 51558 70974 51604
rect 70824 51454 70870 51500
rect 70928 51454 70974 51500
rect 70824 51350 70870 51396
rect 70928 51350 70974 51396
rect 70824 51246 70870 51292
rect 70928 51246 70974 51292
rect 70824 51142 70870 51188
rect 70928 51142 70974 51188
rect 70824 51038 70870 51084
rect 70928 51038 70974 51084
rect 70824 50934 70870 50980
rect 70928 50934 70974 50980
rect 70824 50830 70870 50876
rect 70928 50830 70974 50876
rect 70824 50726 70870 50772
rect 70928 50726 70974 50772
rect 70824 50622 70870 50668
rect 70928 50622 70974 50668
rect 70824 50518 70870 50564
rect 70928 50518 70974 50564
rect 70824 50414 70870 50460
rect 70928 50414 70974 50460
rect 70824 50310 70870 50356
rect 70928 50310 70974 50356
rect 70824 50206 70870 50252
rect 70928 50206 70974 50252
rect 70824 50102 70870 50148
rect 70928 50102 70974 50148
rect 70824 49998 70870 50044
rect 70928 49998 70974 50044
rect 70824 49894 70870 49940
rect 70928 49894 70974 49940
rect 70824 49790 70870 49836
rect 70928 49790 70974 49836
rect 70824 49686 70870 49732
rect 70928 49686 70974 49732
rect 70824 49582 70870 49628
rect 70928 49582 70974 49628
rect 70824 49478 70870 49524
rect 70928 49478 70974 49524
rect 70824 49374 70870 49420
rect 70928 49374 70974 49420
rect 70824 49270 70870 49316
rect 70928 49270 70974 49316
rect 70824 49166 70870 49212
rect 70928 49166 70974 49212
rect 70824 49062 70870 49108
rect 70928 49062 70974 49108
rect 70824 48958 70870 49004
rect 70928 48958 70974 49004
rect 70824 48854 70870 48900
rect 70928 48854 70974 48900
rect 70824 48750 70870 48796
rect 70928 48750 70974 48796
rect 70824 48646 70870 48692
rect 70928 48646 70974 48692
rect 70824 48542 70870 48588
rect 70928 48542 70974 48588
rect 70824 48438 70870 48484
rect 70928 48438 70974 48484
rect 70824 48334 70870 48380
rect 70928 48334 70974 48380
rect 70824 48230 70870 48276
rect 70928 48230 70974 48276
rect 70824 48126 70870 48172
rect 70928 48126 70974 48172
rect 70824 48022 70870 48068
rect 70928 48022 70974 48068
rect 70824 47918 70870 47964
rect 70928 47918 70974 47964
rect 70824 47814 70870 47860
rect 70928 47814 70974 47860
rect 70824 47710 70870 47756
rect 70928 47710 70974 47756
rect 70824 47606 70870 47652
rect 70928 47606 70974 47652
rect 70824 47502 70870 47548
rect 70928 47502 70974 47548
rect 70824 47398 70870 47444
rect 70928 47398 70974 47444
rect 70824 47294 70870 47340
rect 70928 47294 70974 47340
rect 70824 47190 70870 47236
rect 70928 47190 70974 47236
rect 70824 47086 70870 47132
rect 70928 47086 70974 47132
rect 70824 46982 70870 47028
rect 70928 46982 70974 47028
rect 70824 46878 70870 46924
rect 70928 46878 70974 46924
rect 70824 46774 70870 46820
rect 70928 46774 70974 46820
rect 70824 46670 70870 46716
rect 70928 46670 70974 46716
rect 70824 46566 70870 46612
rect 70928 46566 70974 46612
rect 70824 46462 70870 46508
rect 70928 46462 70974 46508
rect 70824 46358 70870 46404
rect 70928 46358 70974 46404
rect 70824 46254 70870 46300
rect 70928 46254 70974 46300
rect 70824 46150 70870 46196
rect 70928 46150 70974 46196
rect 70824 46046 70870 46092
rect 70928 46046 70974 46092
rect 70824 45942 70870 45988
rect 70928 45942 70974 45988
rect 70824 45838 70870 45884
rect 70928 45838 70974 45884
rect 70824 45734 70870 45780
rect 70928 45734 70974 45780
rect 70824 45630 70870 45676
rect 70928 45630 70974 45676
rect 70824 45526 70870 45572
rect 70928 45526 70974 45572
rect 70824 45422 70870 45468
rect 70928 45422 70974 45468
rect 70824 45318 70870 45364
rect 70928 45318 70974 45364
rect 70824 45214 70870 45260
rect 70928 45214 70974 45260
rect 70824 45110 70870 45156
rect 70928 45110 70974 45156
rect 70824 45006 70870 45052
rect 70928 45006 70974 45052
rect 70824 44902 70870 44948
rect 70928 44902 70974 44948
rect 13254 44778 13300 44824
rect 70824 44798 70870 44844
rect 70928 44798 70974 44844
rect 13386 44646 13432 44692
rect 70824 44694 70870 44740
rect 70928 44694 70974 44740
rect 70824 44590 70870 44636
rect 70928 44590 70974 44636
rect 13518 44514 13564 44560
rect 70824 44486 70870 44532
rect 70928 44486 70974 44532
rect 13650 44382 13696 44428
rect 70824 44382 70870 44428
rect 70928 44382 70974 44428
rect 13782 44250 13828 44296
rect 70824 44278 70870 44324
rect 70928 44278 70974 44324
rect 70824 44174 70870 44220
rect 70928 44174 70974 44220
rect 13914 44118 13960 44164
rect 70824 44070 70870 44116
rect 70928 44070 70974 44116
rect 14046 43986 14092 44032
rect 70824 43966 70870 44012
rect 70928 43966 70974 44012
rect 14178 43854 14224 43900
rect 70824 43862 70870 43908
rect 70928 43862 70974 43908
rect 14310 43722 14356 43768
rect 70824 43758 70870 43804
rect 70928 43758 70974 43804
rect 70824 43654 70870 43700
rect 70928 43654 70974 43700
rect 14442 43590 14488 43636
rect 70824 43550 70870 43596
rect 70928 43550 70974 43596
rect 14574 43458 14620 43504
rect 70824 43446 70870 43492
rect 70928 43446 70974 43492
rect 14706 43326 14752 43372
rect 70824 43342 70870 43388
rect 70928 43342 70974 43388
rect 14838 43194 14884 43240
rect 70824 43238 70870 43284
rect 70928 43238 70974 43284
rect 70824 43134 70870 43180
rect 70928 43134 70974 43180
rect 14970 43062 15016 43108
rect 70824 43030 70870 43076
rect 70928 43030 70974 43076
rect 15102 42930 15148 42976
rect 70824 42926 70870 42972
rect 70928 42926 70974 42972
rect 15234 42798 15280 42844
rect 70824 42822 70870 42868
rect 70928 42822 70974 42868
rect 70824 42718 70870 42764
rect 70928 42718 70974 42764
rect 15366 42666 15412 42712
rect 70824 42614 70870 42660
rect 70928 42614 70974 42660
rect 15498 42534 15544 42580
rect 70824 42510 70870 42556
rect 70928 42510 70974 42556
rect 15630 42402 15676 42448
rect 70824 42406 70870 42452
rect 70928 42406 70974 42452
rect 15762 42270 15808 42316
rect 70824 42302 70870 42348
rect 70928 42302 70974 42348
rect 70824 42198 70870 42244
rect 70928 42198 70974 42244
rect 15894 42138 15940 42184
rect 70824 42094 70870 42140
rect 70928 42094 70974 42140
rect 16026 42006 16072 42052
rect 70824 41990 70870 42036
rect 70928 41990 70974 42036
rect 16158 41874 16204 41920
rect 70824 41886 70870 41932
rect 70928 41886 70974 41932
rect 16290 41742 16336 41788
rect 70824 41782 70870 41828
rect 70928 41782 70974 41828
rect 70824 41678 70870 41724
rect 70928 41678 70974 41724
rect 16422 41610 16468 41656
rect 70824 41574 70870 41620
rect 70928 41574 70974 41620
rect 16554 41478 16600 41524
rect 70824 41470 70870 41516
rect 70928 41470 70974 41516
rect 16686 41346 16732 41392
rect 70824 41366 70870 41412
rect 70928 41366 70974 41412
rect 70824 41262 70870 41308
rect 70928 41262 70974 41308
rect 16818 41214 16864 41260
rect 70824 41158 70870 41204
rect 70928 41158 70974 41204
rect 16950 41082 16996 41128
rect 70824 41054 70870 41100
rect 70928 41054 70974 41100
rect 17082 40950 17128 40996
rect 70824 40950 70870 40996
rect 70928 40950 70974 40996
rect 17214 40818 17260 40864
rect 70824 40846 70870 40892
rect 70928 40846 70974 40892
rect 70824 40742 70870 40788
rect 70928 40742 70974 40788
rect 17346 40686 17392 40732
rect 70824 40638 70870 40684
rect 70928 40638 70974 40684
rect 17478 40554 17524 40600
rect 70824 40534 70870 40580
rect 70928 40534 70974 40580
rect 17610 40422 17656 40468
rect 70824 40430 70870 40476
rect 70928 40430 70974 40476
rect 17742 40290 17788 40336
rect 70824 40326 70870 40372
rect 70928 40326 70974 40372
rect 70824 40222 70870 40268
rect 70928 40222 70974 40268
rect 17874 40158 17920 40204
rect 70824 40118 70870 40164
rect 70928 40118 70974 40164
rect 18006 40026 18052 40072
rect 70824 40014 70870 40060
rect 70928 40014 70974 40060
rect 18138 39894 18184 39940
rect 70824 39910 70870 39956
rect 70928 39910 70974 39956
rect 18270 39762 18316 39808
rect 70824 39806 70870 39852
rect 70928 39806 70974 39852
rect 70824 39702 70870 39748
rect 70928 39702 70974 39748
rect 18402 39630 18448 39676
rect 70824 39598 70870 39644
rect 70928 39598 70974 39644
rect 18534 39498 18580 39544
rect 70824 39494 70870 39540
rect 70928 39494 70974 39540
rect 18666 39366 18712 39412
rect 70824 39390 70870 39436
rect 70928 39390 70974 39436
rect 70824 39286 70870 39332
rect 70928 39286 70974 39332
rect 18798 39234 18844 39280
rect 70824 39182 70870 39228
rect 70928 39182 70974 39228
rect 18930 39102 18976 39148
rect 70824 39078 70870 39124
rect 70928 39078 70974 39124
rect 19062 38970 19108 39016
rect 70824 38974 70870 39020
rect 70928 38974 70974 39020
rect 19194 38838 19240 38884
rect 70824 38870 70870 38916
rect 70928 38870 70974 38916
rect 70824 38766 70870 38812
rect 70928 38766 70974 38812
rect 19326 38706 19372 38752
rect 70824 38662 70870 38708
rect 70928 38662 70974 38708
rect 19458 38574 19504 38620
rect 70824 38558 70870 38604
rect 70928 38558 70974 38604
rect 19590 38442 19636 38488
rect 70824 38454 70870 38500
rect 70928 38454 70974 38500
rect 19722 38310 19768 38356
rect 70824 38350 70870 38396
rect 70928 38350 70974 38396
rect 70824 38246 70870 38292
rect 70928 38246 70974 38292
rect 19854 38178 19900 38224
rect 70824 38142 70870 38188
rect 70928 38142 70974 38188
rect 19986 38046 20032 38092
rect 70824 38038 70870 38084
rect 70928 38038 70974 38084
rect 20118 37914 20164 37960
rect 70824 37934 70870 37980
rect 70928 37934 70974 37980
rect 20250 37782 20296 37828
rect 70824 37830 70870 37876
rect 70928 37830 70974 37876
rect 70824 37726 70870 37772
rect 70928 37726 70974 37772
rect 20382 37650 20428 37696
rect 70824 37622 70870 37668
rect 70928 37622 70974 37668
rect 20514 37518 20560 37564
rect 70824 37518 70870 37564
rect 70928 37518 70974 37564
rect 20646 37386 20692 37432
rect 70824 37414 70870 37460
rect 70928 37414 70974 37460
rect 70824 37310 70870 37356
rect 70928 37310 70974 37356
rect 20778 37254 20824 37300
rect 70824 37206 70870 37252
rect 70928 37206 70974 37252
rect 20910 37122 20956 37168
rect 70824 37102 70870 37148
rect 70928 37102 70974 37148
rect 21042 36990 21088 37036
rect 70824 36998 70870 37044
rect 70928 36998 70974 37044
rect 21174 36858 21220 36904
rect 70824 36894 70870 36940
rect 70928 36894 70974 36940
rect 70824 36790 70870 36836
rect 70928 36790 70974 36836
rect 21306 36726 21352 36772
rect 70824 36686 70870 36732
rect 70928 36686 70974 36732
rect 21438 36594 21484 36640
rect 70824 36582 70870 36628
rect 70928 36582 70974 36628
rect 21570 36462 21616 36508
rect 70824 36478 70870 36524
rect 70928 36478 70974 36524
rect 21702 36330 21748 36376
rect 70824 36374 70870 36420
rect 70928 36374 70974 36420
rect 70824 36270 70870 36316
rect 70928 36270 70974 36316
rect 21834 36198 21880 36244
rect 70824 36166 70870 36212
rect 70928 36166 70974 36212
rect 21966 36066 22012 36112
rect 70824 36062 70870 36108
rect 70928 36062 70974 36108
rect 22098 35934 22144 35980
rect 70824 35958 70870 36004
rect 70928 35958 70974 36004
rect 70824 35854 70870 35900
rect 70928 35854 70974 35900
rect 22230 35802 22276 35848
rect 70824 35750 70870 35796
rect 70928 35750 70974 35796
rect 22362 35670 22408 35716
rect 70824 35646 70870 35692
rect 70928 35646 70974 35692
rect 22494 35538 22540 35584
rect 70824 35542 70870 35588
rect 70928 35542 70974 35588
rect 22626 35406 22672 35452
rect 70824 35438 70870 35484
rect 70928 35438 70974 35484
rect 70824 35334 70870 35380
rect 70928 35334 70974 35380
rect 22758 35274 22804 35320
rect 70824 35230 70870 35276
rect 70928 35230 70974 35276
rect 22890 35142 22936 35188
rect 70824 35126 70870 35172
rect 70928 35126 70974 35172
rect 23022 35010 23068 35056
rect 70824 35022 70870 35068
rect 70928 35022 70974 35068
rect 23154 34878 23200 34924
rect 70824 34918 70870 34964
rect 70928 34918 70974 34964
rect 70824 34814 70870 34860
rect 70928 34814 70974 34860
rect 23286 34746 23332 34792
rect 70824 34710 70870 34756
rect 70928 34710 70974 34756
rect 23418 34614 23464 34660
rect 70824 34606 70870 34652
rect 70928 34606 70974 34652
rect 23550 34482 23596 34528
rect 70824 34502 70870 34548
rect 70928 34502 70974 34548
rect 23682 34350 23728 34396
rect 70824 34398 70870 34444
rect 70928 34398 70974 34444
rect 70824 34294 70870 34340
rect 70928 34294 70974 34340
rect 23814 34218 23860 34264
rect 70824 34190 70870 34236
rect 70928 34190 70974 34236
rect 23946 34086 23992 34132
rect 70824 34086 70870 34132
rect 70928 34086 70974 34132
rect 24078 33954 24124 34000
rect 70824 33982 70870 34028
rect 70928 33982 70974 34028
rect 70824 33878 70870 33924
rect 70928 33878 70974 33924
rect 24210 33822 24256 33868
rect 70824 33774 70870 33820
rect 70928 33774 70974 33820
rect 24342 33690 24388 33736
rect 70824 33670 70870 33716
rect 70928 33670 70974 33716
rect 24474 33558 24520 33604
rect 70824 33566 70870 33612
rect 70928 33566 70974 33612
rect 24606 33426 24652 33472
rect 70824 33462 70870 33508
rect 70928 33462 70974 33508
rect 70824 33358 70870 33404
rect 70928 33358 70974 33404
rect 24738 33294 24784 33340
rect 70824 33254 70870 33300
rect 70928 33254 70974 33300
rect 24870 33162 24916 33208
rect 70824 33150 70870 33196
rect 70928 33150 70974 33196
rect 25002 33030 25048 33076
rect 70824 33046 70870 33092
rect 70928 33046 70974 33092
rect 25134 32898 25180 32944
rect 70824 32942 70870 32988
rect 70928 32942 70974 32988
rect 70824 32838 70870 32884
rect 70928 32838 70974 32884
rect 25266 32766 25312 32812
rect 70824 32734 70870 32780
rect 70928 32734 70974 32780
rect 25398 32634 25444 32680
rect 70824 32630 70870 32676
rect 70928 32630 70974 32676
rect 25530 32502 25576 32548
rect 70824 32526 70870 32572
rect 70928 32526 70974 32572
rect 70824 32422 70870 32468
rect 70928 32422 70974 32468
rect 25662 32370 25708 32416
rect 70824 32318 70870 32364
rect 70928 32318 70974 32364
rect 25794 32238 25840 32284
rect 70824 32214 70870 32260
rect 70928 32214 70974 32260
rect 25926 32106 25972 32152
rect 70824 32110 70870 32156
rect 70928 32110 70974 32156
rect 26058 31974 26104 32020
rect 70824 32006 70870 32052
rect 70928 32006 70974 32052
rect 70824 31902 70870 31948
rect 70928 31902 70974 31948
rect 26190 31842 26236 31888
rect 70824 31798 70870 31844
rect 70928 31798 70974 31844
rect 26322 31710 26368 31756
rect 70824 31694 70870 31740
rect 70928 31694 70974 31740
rect 26454 31578 26500 31624
rect 70824 31590 70870 31636
rect 70928 31590 70974 31636
rect 26586 31446 26632 31492
rect 70824 31486 70870 31532
rect 70928 31486 70974 31532
rect 70824 31382 70870 31428
rect 70928 31382 70974 31428
rect 26718 31314 26764 31360
rect 70824 31278 70870 31324
rect 70928 31278 70974 31324
rect 26850 31182 26896 31228
rect 70824 31174 70870 31220
rect 70928 31174 70974 31220
rect 26982 31050 27028 31096
rect 70824 31070 70870 31116
rect 70928 31070 70974 31116
rect 27114 30918 27160 30964
rect 70824 30966 70870 31012
rect 70928 30966 70974 31012
rect 70824 30862 70870 30908
rect 70928 30862 70974 30908
rect 27246 30786 27292 30832
rect 70824 30758 70870 30804
rect 70928 30758 70974 30804
rect 27378 30654 27424 30700
rect 70824 30654 70870 30700
rect 70928 30654 70974 30700
rect 27510 30522 27556 30568
rect 70824 30550 70870 30596
rect 70928 30550 70974 30596
rect 70824 30446 70870 30492
rect 70928 30446 70974 30492
rect 27642 30390 27688 30436
rect 70824 30342 70870 30388
rect 70928 30342 70974 30388
rect 27774 30258 27820 30304
rect 70824 30238 70870 30284
rect 70928 30238 70974 30284
rect 27906 30126 27952 30172
rect 70824 30134 70870 30180
rect 70928 30134 70974 30180
rect 28038 29994 28084 30040
rect 70824 30030 70870 30076
rect 70928 30030 70974 30076
rect 70824 29926 70870 29972
rect 70928 29926 70974 29972
rect 28170 29862 28216 29908
rect 70824 29822 70870 29868
rect 70928 29822 70974 29868
rect 28302 29730 28348 29776
rect 70824 29718 70870 29764
rect 70928 29718 70974 29764
rect 28434 29598 28480 29644
rect 70824 29614 70870 29660
rect 70928 29614 70974 29660
rect 28566 29466 28612 29512
rect 70824 29510 70870 29556
rect 70928 29510 70974 29556
rect 70824 29406 70870 29452
rect 70928 29406 70974 29452
rect 28698 29334 28744 29380
rect 70824 29302 70870 29348
rect 70928 29302 70974 29348
rect 28830 29202 28876 29248
rect 70824 29198 70870 29244
rect 70928 29198 70974 29244
rect 28962 29070 29008 29116
rect 70824 29094 70870 29140
rect 70928 29094 70974 29140
rect 29094 28938 29140 28984
rect 70824 28990 70870 29036
rect 70928 28990 70974 29036
rect 70824 28886 70870 28932
rect 70928 28886 70974 28932
rect 29226 28806 29272 28852
rect 70824 28782 70870 28828
rect 70928 28782 70974 28828
rect 29358 28674 29404 28720
rect 70824 28678 70870 28724
rect 70928 28678 70974 28724
rect 29490 28542 29536 28588
rect 70824 28574 70870 28620
rect 70928 28574 70974 28620
rect 70824 28470 70870 28516
rect 70928 28470 70974 28516
rect 29622 28410 29668 28456
rect 70824 28366 70870 28412
rect 70928 28366 70974 28412
rect 29754 28278 29800 28324
rect 70824 28262 70870 28308
rect 70928 28262 70974 28308
rect 29886 28146 29932 28192
rect 70824 28158 70870 28204
rect 70928 28158 70974 28204
rect 30018 28014 30064 28060
rect 70824 28054 70870 28100
rect 70928 28054 70974 28100
rect 70824 27950 70870 27996
rect 70928 27950 70974 27996
rect 30150 27882 30196 27928
rect 70824 27846 70870 27892
rect 70928 27846 70974 27892
rect 30282 27750 30328 27796
rect 70824 27742 70870 27788
rect 70928 27742 70974 27788
rect 30414 27618 30460 27664
rect 70824 27638 70870 27684
rect 70928 27638 70974 27684
rect 30546 27486 30592 27532
rect 70824 27534 70870 27580
rect 70928 27534 70974 27580
rect 70824 27430 70870 27476
rect 70928 27430 70974 27476
rect 30678 27354 30724 27400
rect 70824 27326 70870 27372
rect 70928 27326 70974 27372
rect 30810 27222 30856 27268
rect 70824 27222 70870 27268
rect 70928 27222 70974 27268
rect 30942 27090 30988 27136
rect 70824 27118 70870 27164
rect 70928 27118 70974 27164
rect 70824 27014 70870 27060
rect 70928 27014 70974 27060
rect 31074 26958 31120 27004
rect 70824 26910 70870 26956
rect 70928 26910 70974 26956
rect 31206 26826 31252 26872
rect 70824 26806 70870 26852
rect 70928 26806 70974 26852
rect 31338 26694 31384 26740
rect 70824 26702 70870 26748
rect 70928 26702 70974 26748
rect 31470 26562 31516 26608
rect 70824 26598 70870 26644
rect 70928 26598 70974 26644
rect 70824 26494 70870 26540
rect 70928 26494 70974 26540
rect 31602 26430 31648 26476
rect 70824 26390 70870 26436
rect 70928 26390 70974 26436
rect 31734 26298 31780 26344
rect 70824 26286 70870 26332
rect 70928 26286 70974 26332
rect 31866 26166 31912 26212
rect 70824 26182 70870 26228
rect 70928 26182 70974 26228
rect 31998 26034 32044 26080
rect 70824 26078 70870 26124
rect 70928 26078 70974 26124
rect 70824 25974 70870 26020
rect 70928 25974 70974 26020
rect 32130 25902 32176 25948
rect 70824 25870 70870 25916
rect 70928 25870 70974 25916
rect 32262 25770 32308 25816
rect 70824 25766 70870 25812
rect 70928 25766 70974 25812
rect 32394 25638 32440 25684
rect 70824 25662 70870 25708
rect 70928 25662 70974 25708
rect 70824 25558 70870 25604
rect 70928 25558 70974 25604
rect 32526 25506 32572 25552
rect 70824 25454 70870 25500
rect 70928 25454 70974 25500
rect 32658 25374 32704 25420
rect 70824 25350 70870 25396
rect 70928 25350 70974 25396
rect 32790 25242 32836 25288
rect 70824 25246 70870 25292
rect 70928 25246 70974 25292
rect 32922 25110 32968 25156
rect 70824 25142 70870 25188
rect 70928 25142 70974 25188
rect 70824 25038 70870 25084
rect 70928 25038 70974 25084
rect 33054 24978 33100 25024
rect 70824 24934 70870 24980
rect 70928 24934 70974 24980
rect 33186 24846 33232 24892
rect 70824 24830 70870 24876
rect 70928 24830 70974 24876
rect 33318 24714 33364 24760
rect 70824 24726 70870 24772
rect 70928 24726 70974 24772
rect 33450 24582 33496 24628
rect 70824 24622 70870 24668
rect 70928 24622 70974 24668
rect 70824 24518 70870 24564
rect 70928 24518 70974 24564
rect 33582 24450 33628 24496
rect 70824 24414 70870 24460
rect 70928 24414 70974 24460
rect 33714 24318 33760 24364
rect 70824 24310 70870 24356
rect 70928 24310 70974 24356
rect 33846 24186 33892 24232
rect 70824 24206 70870 24252
rect 70928 24206 70974 24252
rect 33978 24054 34024 24100
rect 70824 24102 70870 24148
rect 70928 24102 70974 24148
rect 70824 23998 70870 24044
rect 70928 23998 70974 24044
rect 34110 23922 34156 23968
rect 70824 23894 70870 23940
rect 70928 23894 70974 23940
rect 34242 23790 34288 23836
rect 70824 23790 70870 23836
rect 70928 23790 70974 23836
rect 34374 23658 34420 23704
rect 70824 23686 70870 23732
rect 70928 23686 70974 23732
rect 70824 23582 70870 23628
rect 70928 23582 70974 23628
rect 34506 23526 34552 23572
rect 70824 23478 70870 23524
rect 70928 23478 70974 23524
rect 34638 23394 34684 23440
rect 70824 23374 70870 23420
rect 70928 23374 70974 23420
rect 34770 23262 34816 23308
rect 70824 23270 70870 23316
rect 70928 23270 70974 23316
rect 34902 23130 34948 23176
rect 70824 23166 70870 23212
rect 70928 23166 70974 23212
rect 70824 23062 70870 23108
rect 70928 23062 70974 23108
rect 35034 22998 35080 23044
rect 70824 22958 70870 23004
rect 70928 22958 70974 23004
rect 35166 22866 35212 22912
rect 70824 22854 70870 22900
rect 70928 22854 70974 22900
rect 35298 22734 35344 22780
rect 70824 22750 70870 22796
rect 70928 22750 70974 22796
rect 35430 22602 35476 22648
rect 70824 22646 70870 22692
rect 70928 22646 70974 22692
rect 70824 22542 70870 22588
rect 70928 22542 70974 22588
rect 35562 22470 35608 22516
rect 70824 22438 70870 22484
rect 70928 22438 70974 22484
rect 35694 22338 35740 22384
rect 70824 22334 70870 22380
rect 70928 22334 70974 22380
rect 35826 22206 35872 22252
rect 70824 22230 70870 22276
rect 70928 22230 70974 22276
rect 70824 22126 70870 22172
rect 70928 22126 70974 22172
rect 35958 22074 36004 22120
rect 70824 22022 70870 22068
rect 70928 22022 70974 22068
rect 36090 21942 36136 21988
rect 70824 21918 70870 21964
rect 70928 21918 70974 21964
rect 36222 21810 36268 21856
rect 70824 21814 70870 21860
rect 70928 21814 70974 21860
rect 36354 21678 36400 21724
rect 70824 21710 70870 21756
rect 70928 21710 70974 21756
rect 70824 21606 70870 21652
rect 70928 21606 70974 21652
rect 36486 21546 36532 21592
rect 70824 21502 70870 21548
rect 70928 21502 70974 21548
rect 36618 21414 36664 21460
rect 70824 21398 70870 21444
rect 70928 21398 70974 21444
rect 36750 21282 36796 21328
rect 70824 21294 70870 21340
rect 70928 21294 70974 21340
rect 36882 21150 36928 21196
rect 70824 21190 70870 21236
rect 70928 21190 70974 21236
rect 70824 21086 70870 21132
rect 70928 21086 70974 21132
rect 37014 21018 37060 21064
rect 70824 20982 70870 21028
rect 70928 20982 70974 21028
rect 37146 20886 37192 20932
rect 70824 20878 70870 20924
rect 70928 20878 70974 20924
rect 37278 20754 37324 20800
rect 70824 20774 70870 20820
rect 70928 20774 70974 20820
rect 37410 20622 37456 20668
rect 70824 20670 70870 20716
rect 70928 20670 70974 20716
rect 70824 20566 70870 20612
rect 70928 20566 70974 20612
rect 37542 20490 37588 20536
rect 70824 20462 70870 20508
rect 70928 20462 70974 20508
rect 37674 20358 37720 20404
rect 70824 20358 70870 20404
rect 70928 20358 70974 20404
rect 37806 20226 37852 20272
rect 70824 20254 70870 20300
rect 70928 20254 70974 20300
rect 70824 20150 70870 20196
rect 70928 20150 70974 20196
rect 37938 20094 37984 20140
rect 70824 20046 70870 20092
rect 70928 20046 70974 20092
rect 38070 19962 38116 20008
rect 70824 19942 70870 19988
rect 70928 19942 70974 19988
rect 38202 19830 38248 19876
rect 70824 19838 70870 19884
rect 70928 19838 70974 19884
rect 38334 19698 38380 19744
rect 70824 19734 70870 19780
rect 70928 19734 70974 19780
rect 70824 19630 70870 19676
rect 70928 19630 70974 19676
rect 38466 19566 38512 19612
rect 70824 19526 70870 19572
rect 70928 19526 70974 19572
rect 38598 19434 38644 19480
rect 70824 19422 70870 19468
rect 70928 19422 70974 19468
rect 38730 19302 38776 19348
rect 70824 19318 70870 19364
rect 70928 19318 70974 19364
rect 38862 19170 38908 19216
rect 70824 19214 70870 19260
rect 70928 19214 70974 19260
rect 70824 19110 70870 19156
rect 70928 19110 70974 19156
rect 38994 19038 39040 19084
rect 70824 19006 70870 19052
rect 70928 19006 70974 19052
rect 39126 18906 39172 18952
rect 70824 18902 70870 18948
rect 70928 18902 70974 18948
rect 39258 18774 39304 18820
rect 70824 18798 70870 18844
rect 70928 18798 70974 18844
rect 70824 18694 70870 18740
rect 70928 18694 70974 18740
rect 39390 18642 39436 18688
rect 70824 18590 70870 18636
rect 70928 18590 70974 18636
rect 39522 18510 39568 18556
rect 70824 18486 70870 18532
rect 70928 18486 70974 18532
rect 39654 18378 39700 18424
rect 70824 18382 70870 18428
rect 70928 18382 70974 18428
rect 39786 18246 39832 18292
rect 70824 18278 70870 18324
rect 70928 18278 70974 18324
rect 70824 18174 70870 18220
rect 70928 18174 70974 18220
rect 39918 18114 39964 18160
rect 70824 18070 70870 18116
rect 70928 18070 70974 18116
rect 40050 17982 40096 18028
rect 70824 17966 70870 18012
rect 70928 17966 70974 18012
rect 40182 17850 40228 17896
rect 70824 17862 70870 17908
rect 70928 17862 70974 17908
rect 40314 17718 40360 17764
rect 70824 17758 70870 17804
rect 70928 17758 70974 17804
rect 70824 17654 70870 17700
rect 70928 17654 70974 17700
rect 40446 17586 40492 17632
rect 70824 17550 70870 17596
rect 70928 17550 70974 17596
rect 40578 17454 40624 17500
rect 70824 17446 70870 17492
rect 70928 17446 70974 17492
rect 40710 17322 40756 17368
rect 70824 17342 70870 17388
rect 70928 17342 70974 17388
rect 70824 17238 70870 17284
rect 70928 17238 70974 17284
rect 40842 17190 40888 17236
rect 70824 17134 70870 17180
rect 70928 17134 70974 17180
rect 40974 17058 41020 17104
rect 70824 17030 70870 17076
rect 70928 17030 70974 17076
rect 41106 16926 41152 16972
rect 70824 16926 70870 16972
rect 70928 16926 70974 16972
rect 41238 16794 41284 16840
rect 70824 16822 70870 16868
rect 70928 16822 70974 16868
rect 70824 16718 70870 16764
rect 70928 16718 70974 16764
rect 41370 16662 41416 16708
rect 70824 16614 70870 16660
rect 70928 16614 70974 16660
rect 41502 16530 41548 16576
rect 70824 16510 70870 16556
rect 70928 16510 70974 16556
rect 41634 16398 41680 16444
rect 70824 16406 70870 16452
rect 70928 16406 70974 16452
rect 41766 16266 41812 16312
rect 70824 16302 70870 16348
rect 70928 16302 70974 16348
rect 70824 16198 70870 16244
rect 70928 16198 70974 16244
rect 41898 16134 41944 16180
rect 70824 16094 70870 16140
rect 70928 16094 70974 16140
rect 42030 16002 42076 16048
rect 70824 15990 70870 16036
rect 70928 15990 70974 16036
rect 42162 15870 42208 15916
rect 70824 15886 70870 15932
rect 70928 15886 70974 15932
rect 42294 15738 42340 15784
rect 70824 15782 70870 15828
rect 70928 15782 70974 15828
rect 70824 15678 70870 15724
rect 70928 15678 70974 15724
rect 42426 15606 42472 15652
rect 70824 15574 70870 15620
rect 70928 15574 70974 15620
rect 42558 15474 42604 15520
rect 70824 15470 70870 15516
rect 70928 15470 70974 15516
rect 42690 15342 42736 15388
rect 70824 15366 70870 15412
rect 70928 15366 70974 15412
rect 70824 15262 70870 15308
rect 70928 15262 70974 15308
rect 42822 15210 42868 15256
rect 70824 15158 70870 15204
rect 70928 15158 70974 15204
rect 42954 15078 43000 15124
rect 70824 15054 70870 15100
rect 70928 15054 70974 15100
rect 43086 14946 43132 14992
rect 70824 14950 70870 14996
rect 70928 14950 70974 14996
rect 43218 14814 43264 14860
rect 70824 14846 70870 14892
rect 70928 14846 70974 14892
rect 70824 14742 70870 14788
rect 70928 14742 70974 14788
rect 43350 14682 43396 14728
rect 70824 14638 70870 14684
rect 70928 14638 70974 14684
rect 43482 14550 43528 14596
rect 70824 14534 70870 14580
rect 70928 14534 70974 14580
rect 43614 14418 43660 14464
rect 70824 14430 70870 14476
rect 70928 14430 70974 14476
rect 43746 14286 43792 14332
rect 70824 14326 70870 14372
rect 70928 14326 70974 14372
rect 70824 14222 70870 14268
rect 70928 14222 70974 14268
rect 43878 14154 43924 14200
rect 70824 14118 70870 14164
rect 70928 14118 70974 14164
rect 44010 14022 44056 14068
rect 70824 14014 70870 14060
rect 70928 14014 70974 14060
rect 44142 13890 44188 13936
rect 70824 13910 70870 13956
rect 70928 13910 70974 13956
rect 44274 13758 44320 13804
rect 70824 13806 70870 13852
rect 70928 13806 70974 13852
rect 70824 13702 70870 13748
rect 70928 13702 70974 13748
rect 44406 13626 44452 13672
rect 70824 13598 70870 13644
rect 70928 13598 70974 13644
rect 44538 13494 44584 13540
rect 70824 13494 70870 13540
rect 70928 13494 70974 13540
rect 44670 13362 44716 13408
rect 70824 13390 70870 13436
rect 70928 13390 70974 13436
rect 44850 13210 44896 13256
rect 45088 13223 45134 13269
rect 45192 13223 45238 13269
rect 45296 13223 45342 13269
rect 45400 13223 45446 13269
rect 45504 13223 45550 13269
rect 45608 13223 45654 13269
rect 45712 13223 45758 13269
rect 45816 13223 45862 13269
rect 45920 13223 45966 13269
rect 46024 13223 46070 13269
rect 46128 13223 46174 13269
rect 46232 13223 46278 13269
rect 46336 13223 46382 13269
rect 46440 13223 46486 13269
rect 46544 13223 46590 13269
rect 46648 13223 46694 13269
rect 46752 13223 46798 13269
rect 46856 13223 46902 13269
rect 46960 13223 47006 13269
rect 47064 13223 47110 13269
rect 47168 13223 47214 13269
rect 47272 13223 47318 13269
rect 47376 13223 47422 13269
rect 47480 13223 47526 13269
rect 47584 13223 47630 13269
rect 47688 13223 47734 13269
rect 47792 13223 47838 13269
rect 47896 13223 47942 13269
rect 48000 13223 48046 13269
rect 48104 13223 48150 13269
rect 48208 13223 48254 13269
rect 48312 13223 48358 13269
rect 48416 13223 48462 13269
rect 48520 13223 48566 13269
rect 48624 13223 48670 13269
rect 48728 13223 48774 13269
rect 48832 13223 48878 13269
rect 48936 13223 48982 13269
rect 49040 13223 49086 13269
rect 49144 13223 49190 13269
rect 49248 13223 49294 13269
rect 49352 13223 49398 13269
rect 49456 13223 49502 13269
rect 49560 13223 49606 13269
rect 49664 13223 49710 13269
rect 49768 13223 49814 13269
rect 49872 13223 49918 13269
rect 49976 13223 50022 13269
rect 50080 13223 50126 13269
rect 50184 13223 50230 13269
rect 50288 13223 50334 13269
rect 50392 13223 50438 13269
rect 50496 13223 50542 13269
rect 50600 13223 50646 13269
rect 50704 13223 50750 13269
rect 50808 13223 50854 13269
rect 50912 13223 50958 13269
rect 51016 13223 51062 13269
rect 51120 13223 51166 13269
rect 51224 13223 51270 13269
rect 51328 13223 51374 13269
rect 51432 13223 51478 13269
rect 51536 13223 51582 13269
rect 51640 13223 51686 13269
rect 51744 13223 51790 13269
rect 51848 13223 51894 13269
rect 51952 13223 51998 13269
rect 52056 13223 52102 13269
rect 52160 13223 52206 13269
rect 52264 13223 52310 13269
rect 52368 13223 52414 13269
rect 52472 13223 52518 13269
rect 52576 13223 52622 13269
rect 52680 13223 52726 13269
rect 52784 13223 52830 13269
rect 52888 13223 52934 13269
rect 52992 13223 53038 13269
rect 53096 13223 53142 13269
rect 53200 13223 53246 13269
rect 53304 13223 53350 13269
rect 53408 13223 53454 13269
rect 53512 13223 53558 13269
rect 53616 13223 53662 13269
rect 53720 13223 53766 13269
rect 53824 13223 53870 13269
rect 53928 13223 53974 13269
rect 54032 13223 54078 13269
rect 54136 13223 54182 13269
rect 54240 13223 54286 13269
rect 54344 13223 54390 13269
rect 54448 13223 54494 13269
rect 54552 13223 54598 13269
rect 54656 13223 54702 13269
rect 54760 13223 54806 13269
rect 54864 13223 54910 13269
rect 54968 13223 55014 13269
rect 55072 13223 55118 13269
rect 55176 13223 55222 13269
rect 55280 13223 55326 13269
rect 55384 13223 55430 13269
rect 55488 13223 55534 13269
rect 55592 13223 55638 13269
rect 55696 13223 55742 13269
rect 55800 13223 55846 13269
rect 55904 13223 55950 13269
rect 56008 13223 56054 13269
rect 56112 13223 56158 13269
rect 56216 13223 56262 13269
rect 56320 13223 56366 13269
rect 56424 13223 56470 13269
rect 56528 13223 56574 13269
rect 56632 13223 56678 13269
rect 56736 13223 56782 13269
rect 56840 13223 56886 13269
rect 56944 13223 56990 13269
rect 57048 13223 57094 13269
rect 57152 13223 57198 13269
rect 57256 13223 57302 13269
rect 57360 13223 57406 13269
rect 57464 13223 57510 13269
rect 57568 13223 57614 13269
rect 57672 13223 57718 13269
rect 57776 13223 57822 13269
rect 57880 13223 57926 13269
rect 57984 13223 58030 13269
rect 58088 13223 58134 13269
rect 58192 13223 58238 13269
rect 58296 13223 58342 13269
rect 58400 13223 58446 13269
rect 58504 13223 58550 13269
rect 58608 13223 58654 13269
rect 58712 13223 58758 13269
rect 58816 13223 58862 13269
rect 58920 13223 58966 13269
rect 59024 13223 59070 13269
rect 59128 13223 59174 13269
rect 59232 13223 59278 13269
rect 59336 13223 59382 13269
rect 59440 13223 59486 13269
rect 59544 13223 59590 13269
rect 59648 13223 59694 13269
rect 59752 13223 59798 13269
rect 59856 13223 59902 13269
rect 59960 13223 60006 13269
rect 60064 13223 60110 13269
rect 60168 13223 60214 13269
rect 60272 13223 60318 13269
rect 60376 13223 60422 13269
rect 60480 13223 60526 13269
rect 60584 13223 60630 13269
rect 60688 13223 60734 13269
rect 60792 13223 60838 13269
rect 60896 13223 60942 13269
rect 61000 13223 61046 13269
rect 61104 13223 61150 13269
rect 61208 13223 61254 13269
rect 61312 13223 61358 13269
rect 61416 13223 61462 13269
rect 61520 13223 61566 13269
rect 61624 13223 61670 13269
rect 61728 13223 61774 13269
rect 61832 13223 61878 13269
rect 61936 13223 61982 13269
rect 62040 13223 62086 13269
rect 62144 13223 62190 13269
rect 62248 13223 62294 13269
rect 62352 13223 62398 13269
rect 62456 13223 62502 13269
rect 62560 13223 62606 13269
rect 62664 13223 62710 13269
rect 62768 13223 62814 13269
rect 62872 13223 62918 13269
rect 62976 13223 63022 13269
rect 63080 13223 63126 13269
rect 63184 13223 63230 13269
rect 63288 13223 63334 13269
rect 63392 13223 63438 13269
rect 63496 13223 63542 13269
rect 63600 13223 63646 13269
rect 63704 13223 63750 13269
rect 63808 13223 63854 13269
rect 63912 13223 63958 13269
rect 64016 13223 64062 13269
rect 64120 13223 64166 13269
rect 64224 13223 64270 13269
rect 64328 13223 64374 13269
rect 64432 13223 64478 13269
rect 64536 13223 64582 13269
rect 64640 13223 64686 13269
rect 64744 13223 64790 13269
rect 64848 13223 64894 13269
rect 64952 13223 64998 13269
rect 65056 13223 65102 13269
rect 65160 13223 65206 13269
rect 65264 13223 65310 13269
rect 65368 13223 65414 13269
rect 65472 13223 65518 13269
rect 65576 13223 65622 13269
rect 65680 13223 65726 13269
rect 65784 13223 65830 13269
rect 65888 13223 65934 13269
rect 65992 13223 66038 13269
rect 66096 13223 66142 13269
rect 66200 13223 66246 13269
rect 66304 13223 66350 13269
rect 66408 13223 66454 13269
rect 66512 13223 66558 13269
rect 66616 13223 66662 13269
rect 66720 13223 66766 13269
rect 66824 13223 66870 13269
rect 66928 13223 66974 13269
rect 67032 13223 67078 13269
rect 67136 13223 67182 13269
rect 67240 13223 67286 13269
rect 67344 13223 67390 13269
rect 67448 13223 67494 13269
rect 67552 13223 67598 13269
rect 67656 13223 67702 13269
rect 67760 13223 67806 13269
rect 67864 13223 67910 13269
rect 67968 13223 68014 13269
rect 68072 13223 68118 13269
rect 68176 13223 68222 13269
rect 68280 13223 68326 13269
rect 68384 13223 68430 13269
rect 68488 13223 68534 13269
rect 68592 13223 68638 13269
rect 68696 13223 68742 13269
rect 68800 13223 68846 13269
rect 68904 13223 68950 13269
rect 69008 13223 69054 13269
rect 69112 13223 69158 13269
rect 69216 13223 69262 13269
rect 69320 13223 69366 13269
rect 69424 13223 69470 13269
rect 69528 13223 69574 13269
rect 69632 13223 69678 13269
rect 69736 13223 69782 13269
rect 69840 13223 69886 13269
rect 69944 13223 69990 13269
rect 70048 13223 70094 13269
rect 70152 13223 70198 13269
rect 70256 13223 70302 13269
rect 70360 13223 70406 13269
rect 70464 13223 70510 13269
rect 70568 13223 70614 13269
rect 70672 13223 70718 13269
rect 70776 13223 70822 13269
rect 70880 13223 70926 13269
rect 45088 13119 45134 13165
rect 45192 13119 45238 13165
rect 45296 13119 45342 13165
rect 45400 13119 45446 13165
rect 45504 13119 45550 13165
rect 45608 13119 45654 13165
rect 45712 13119 45758 13165
rect 45816 13119 45862 13165
rect 45920 13119 45966 13165
rect 46024 13119 46070 13165
rect 46128 13119 46174 13165
rect 46232 13119 46278 13165
rect 46336 13119 46382 13165
rect 46440 13119 46486 13165
rect 46544 13119 46590 13165
rect 46648 13119 46694 13165
rect 46752 13119 46798 13165
rect 46856 13119 46902 13165
rect 46960 13119 47006 13165
rect 47064 13119 47110 13165
rect 47168 13119 47214 13165
rect 47272 13119 47318 13165
rect 47376 13119 47422 13165
rect 47480 13119 47526 13165
rect 47584 13119 47630 13165
rect 47688 13119 47734 13165
rect 47792 13119 47838 13165
rect 47896 13119 47942 13165
rect 48000 13119 48046 13165
rect 48104 13119 48150 13165
rect 48208 13119 48254 13165
rect 48312 13119 48358 13165
rect 48416 13119 48462 13165
rect 48520 13119 48566 13165
rect 48624 13119 48670 13165
rect 48728 13119 48774 13165
rect 48832 13119 48878 13165
rect 48936 13119 48982 13165
rect 49040 13119 49086 13165
rect 49144 13119 49190 13165
rect 49248 13119 49294 13165
rect 49352 13119 49398 13165
rect 49456 13119 49502 13165
rect 49560 13119 49606 13165
rect 49664 13119 49710 13165
rect 49768 13119 49814 13165
rect 49872 13119 49918 13165
rect 49976 13119 50022 13165
rect 50080 13119 50126 13165
rect 50184 13119 50230 13165
rect 50288 13119 50334 13165
rect 50392 13119 50438 13165
rect 50496 13119 50542 13165
rect 50600 13119 50646 13165
rect 50704 13119 50750 13165
rect 50808 13119 50854 13165
rect 50912 13119 50958 13165
rect 51016 13119 51062 13165
rect 51120 13119 51166 13165
rect 51224 13119 51270 13165
rect 51328 13119 51374 13165
rect 51432 13119 51478 13165
rect 51536 13119 51582 13165
rect 51640 13119 51686 13165
rect 51744 13119 51790 13165
rect 51848 13119 51894 13165
rect 51952 13119 51998 13165
rect 52056 13119 52102 13165
rect 52160 13119 52206 13165
rect 52264 13119 52310 13165
rect 52368 13119 52414 13165
rect 52472 13119 52518 13165
rect 52576 13119 52622 13165
rect 52680 13119 52726 13165
rect 52784 13119 52830 13165
rect 52888 13119 52934 13165
rect 52992 13119 53038 13165
rect 53096 13119 53142 13165
rect 53200 13119 53246 13165
rect 53304 13119 53350 13165
rect 53408 13119 53454 13165
rect 53512 13119 53558 13165
rect 53616 13119 53662 13165
rect 53720 13119 53766 13165
rect 53824 13119 53870 13165
rect 53928 13119 53974 13165
rect 54032 13119 54078 13165
rect 54136 13119 54182 13165
rect 54240 13119 54286 13165
rect 54344 13119 54390 13165
rect 54448 13119 54494 13165
rect 54552 13119 54598 13165
rect 54656 13119 54702 13165
rect 54760 13119 54806 13165
rect 54864 13119 54910 13165
rect 54968 13119 55014 13165
rect 55072 13119 55118 13165
rect 55176 13119 55222 13165
rect 55280 13119 55326 13165
rect 55384 13119 55430 13165
rect 55488 13119 55534 13165
rect 55592 13119 55638 13165
rect 55696 13119 55742 13165
rect 55800 13119 55846 13165
rect 55904 13119 55950 13165
rect 56008 13119 56054 13165
rect 56112 13119 56158 13165
rect 56216 13119 56262 13165
rect 56320 13119 56366 13165
rect 56424 13119 56470 13165
rect 56528 13119 56574 13165
rect 56632 13119 56678 13165
rect 56736 13119 56782 13165
rect 56840 13119 56886 13165
rect 56944 13119 56990 13165
rect 57048 13119 57094 13165
rect 57152 13119 57198 13165
rect 57256 13119 57302 13165
rect 57360 13119 57406 13165
rect 57464 13119 57510 13165
rect 57568 13119 57614 13165
rect 57672 13119 57718 13165
rect 57776 13119 57822 13165
rect 57880 13119 57926 13165
rect 57984 13119 58030 13165
rect 58088 13119 58134 13165
rect 58192 13119 58238 13165
rect 58296 13119 58342 13165
rect 58400 13119 58446 13165
rect 58504 13119 58550 13165
rect 58608 13119 58654 13165
rect 58712 13119 58758 13165
rect 58816 13119 58862 13165
rect 58920 13119 58966 13165
rect 59024 13119 59070 13165
rect 59128 13119 59174 13165
rect 59232 13119 59278 13165
rect 59336 13119 59382 13165
rect 59440 13119 59486 13165
rect 59544 13119 59590 13165
rect 59648 13119 59694 13165
rect 59752 13119 59798 13165
rect 59856 13119 59902 13165
rect 59960 13119 60006 13165
rect 60064 13119 60110 13165
rect 60168 13119 60214 13165
rect 60272 13119 60318 13165
rect 60376 13119 60422 13165
rect 60480 13119 60526 13165
rect 60584 13119 60630 13165
rect 60688 13119 60734 13165
rect 60792 13119 60838 13165
rect 60896 13119 60942 13165
rect 61000 13119 61046 13165
rect 61104 13119 61150 13165
rect 61208 13119 61254 13165
rect 61312 13119 61358 13165
rect 61416 13119 61462 13165
rect 61520 13119 61566 13165
rect 61624 13119 61670 13165
rect 61728 13119 61774 13165
rect 61832 13119 61878 13165
rect 61936 13119 61982 13165
rect 62040 13119 62086 13165
rect 62144 13119 62190 13165
rect 62248 13119 62294 13165
rect 62352 13119 62398 13165
rect 62456 13119 62502 13165
rect 62560 13119 62606 13165
rect 62664 13119 62710 13165
rect 62768 13119 62814 13165
rect 62872 13119 62918 13165
rect 62976 13119 63022 13165
rect 63080 13119 63126 13165
rect 63184 13119 63230 13165
rect 63288 13119 63334 13165
rect 63392 13119 63438 13165
rect 63496 13119 63542 13165
rect 63600 13119 63646 13165
rect 63704 13119 63750 13165
rect 63808 13119 63854 13165
rect 63912 13119 63958 13165
rect 64016 13119 64062 13165
rect 64120 13119 64166 13165
rect 64224 13119 64270 13165
rect 64328 13119 64374 13165
rect 64432 13119 64478 13165
rect 64536 13119 64582 13165
rect 64640 13119 64686 13165
rect 64744 13119 64790 13165
rect 64848 13119 64894 13165
rect 64952 13119 64998 13165
rect 65056 13119 65102 13165
rect 65160 13119 65206 13165
rect 65264 13119 65310 13165
rect 65368 13119 65414 13165
rect 65472 13119 65518 13165
rect 65576 13119 65622 13165
rect 65680 13119 65726 13165
rect 65784 13119 65830 13165
rect 65888 13119 65934 13165
rect 65992 13119 66038 13165
rect 66096 13119 66142 13165
rect 66200 13119 66246 13165
rect 66304 13119 66350 13165
rect 66408 13119 66454 13165
rect 66512 13119 66558 13165
rect 66616 13119 66662 13165
rect 66720 13119 66766 13165
rect 66824 13119 66870 13165
rect 66928 13119 66974 13165
rect 67032 13119 67078 13165
rect 67136 13119 67182 13165
rect 67240 13119 67286 13165
rect 67344 13119 67390 13165
rect 67448 13119 67494 13165
rect 67552 13119 67598 13165
rect 67656 13119 67702 13165
rect 67760 13119 67806 13165
rect 67864 13119 67910 13165
rect 67968 13119 68014 13165
rect 68072 13119 68118 13165
rect 68176 13119 68222 13165
rect 68280 13119 68326 13165
rect 68384 13119 68430 13165
rect 68488 13119 68534 13165
rect 68592 13119 68638 13165
rect 68696 13119 68742 13165
rect 68800 13119 68846 13165
rect 68904 13119 68950 13165
rect 69008 13119 69054 13165
rect 69112 13119 69158 13165
rect 69216 13119 69262 13165
rect 69320 13119 69366 13165
rect 69424 13119 69470 13165
rect 69528 13119 69574 13165
rect 69632 13119 69678 13165
rect 69736 13119 69782 13165
rect 69840 13119 69886 13165
rect 69944 13119 69990 13165
rect 70048 13119 70094 13165
rect 70152 13119 70198 13165
rect 70256 13119 70302 13165
rect 70360 13119 70406 13165
rect 70464 13119 70510 13165
rect 70568 13119 70614 13165
rect 70672 13119 70718 13165
rect 70776 13119 70822 13165
rect 70880 13119 70926 13165
<< metal1 >>
rect 13108 70975 69957 71000
rect 13108 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69957 70975
rect 13108 70871 69957 70929
rect 13108 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69957 70871
rect 13108 70814 69957 70825
rect 13108 70767 13280 70814
rect 13108 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13280 70767
rect 13108 70663 13280 70721
rect 13108 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13280 70663
rect 13108 70559 13280 70617
rect 13108 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13280 70559
rect 13108 70455 13280 70513
rect 13108 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13280 70455
rect 13108 70351 13280 70409
rect 13108 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13280 70351
rect 13108 70247 13280 70305
rect 13108 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13280 70247
rect 13108 70143 13280 70201
rect 13108 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13280 70143
rect 13108 70039 13280 70097
rect 13108 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13280 70039
rect 13108 69935 13280 69993
rect 13108 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13280 69935
rect 13108 69831 13280 69889
rect 13108 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13280 69831
rect 69785 70720 69957 70814
rect 69785 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69957 70720
rect 69785 70616 69957 70674
rect 69785 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69957 70616
rect 69785 70512 69957 70570
rect 69785 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69957 70512
rect 69785 70408 69957 70466
rect 69785 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69957 70408
rect 69785 70304 69957 70362
rect 69785 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69957 70304
rect 69785 70200 69957 70258
rect 69785 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69957 70200
rect 69785 70096 69957 70154
rect 69785 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69957 70096
rect 69785 69957 69957 70050
rect 69785 69946 71000 69957
rect 69785 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69785 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69785 69842 71000 69862
rect 69785 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69785 69785 70824 69796
rect 13108 69727 13280 69785
rect 13108 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13280 69727
rect 13108 69623 13280 69681
rect 13108 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13280 69623
rect 13108 69519 13280 69577
rect 13108 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13280 69519
rect 13108 69415 13280 69473
rect 13108 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13280 69415
rect 13108 69311 13280 69369
rect 13108 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13280 69311
rect 13108 69207 13280 69265
rect 13108 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13280 69207
rect 13108 69103 13280 69161
rect 13108 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13280 69103
rect 13108 68999 13280 69057
rect 13108 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13280 68999
rect 13108 68895 13280 68953
rect 13108 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13280 68895
rect 13108 68791 13280 68849
rect 13108 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13280 68791
rect 13108 68687 13280 68745
rect 13108 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13280 68687
rect 13108 68583 13280 68641
rect 13108 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13280 68583
rect 13108 68479 13280 68537
rect 13108 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13280 68479
rect 13108 68375 13280 68433
rect 13108 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13280 68375
rect 13108 68271 13280 68329
rect 13108 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13280 68271
rect 13108 68167 13280 68225
rect 13108 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13280 68167
rect 13108 68063 13280 68121
rect 13108 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13280 68063
rect 13108 67959 13280 68017
rect 13108 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13280 67959
rect 13108 67855 13280 67913
rect 13108 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13280 67855
rect 13108 67751 13280 67809
rect 13108 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13280 67751
rect 13108 67647 13280 67705
rect 13108 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13280 67647
rect 13108 67543 13280 67601
rect 13108 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13280 67543
rect 13108 67439 13280 67497
rect 13108 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13280 67439
rect 13108 67335 13280 67393
rect 13108 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13280 67335
rect 13108 67231 13280 67289
rect 13108 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13280 67231
rect 13108 67127 13280 67185
rect 13108 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13280 67127
rect 13108 67023 13280 67081
rect 13108 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13280 67023
rect 13108 66919 13280 66977
rect 13108 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13280 66919
rect 13108 66815 13280 66873
rect 13108 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13280 66815
rect 13108 66711 13280 66769
rect 13108 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13280 66711
rect 13108 66607 13280 66665
rect 13108 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13280 66607
rect 13108 66503 13280 66561
rect 13108 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13280 66503
rect 13108 66399 13280 66457
rect 13108 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13280 66399
rect 13108 66295 13280 66353
rect 13108 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13280 66295
rect 13108 66191 13280 66249
rect 13108 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13280 66191
rect 13108 66087 13280 66145
rect 13108 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13280 66087
rect 13108 65983 13280 66041
rect 13108 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13280 65983
rect 13108 65879 13280 65937
rect 13108 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13280 65879
rect 13108 65775 13280 65833
rect 13108 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13280 65775
rect 13108 65671 13280 65729
rect 13108 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13280 65671
rect 13108 65567 13280 65625
rect 13108 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13280 65567
rect 13108 65463 13280 65521
rect 13108 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13280 65463
rect 13108 65359 13280 65417
rect 13108 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13280 65359
rect 13108 65255 13280 65313
rect 13108 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13280 65255
rect 13108 65151 13280 65209
rect 13108 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13280 65151
rect 13108 65047 13280 65105
rect 13108 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13280 65047
rect 13108 64943 13280 65001
rect 13108 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13280 64943
rect 13108 64839 13280 64897
rect 13108 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13280 64839
rect 13108 64735 13280 64793
rect 13108 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13280 64735
rect 13108 64631 13280 64689
rect 13108 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13280 64631
rect 13108 64527 13280 64585
rect 13108 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13280 64527
rect 13108 64423 13280 64481
rect 13108 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13280 64423
rect 13108 64319 13280 64377
rect 13108 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13280 64319
rect 13108 64215 13280 64273
rect 13108 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13280 64215
rect 13108 64111 13280 64169
rect 13108 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13280 64111
rect 13108 64007 13280 64065
rect 13108 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13280 64007
rect 13108 63903 13280 63961
rect 13108 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13280 63903
rect 13108 63799 13280 63857
rect 13108 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13280 63799
rect 13108 63695 13280 63753
rect 13108 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13280 63695
rect 13108 63591 13280 63649
rect 13108 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13280 63591
rect 13108 63487 13280 63545
rect 13108 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13280 63487
rect 13108 63383 13280 63441
rect 13108 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13280 63383
rect 13108 63279 13280 63337
rect 13108 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13280 63279
rect 13108 63175 13280 63233
rect 13108 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13280 63175
rect 13108 63071 13280 63129
rect 13108 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13280 63071
rect 13108 62967 13280 63025
rect 13108 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13280 62967
rect 13108 62863 13280 62921
rect 13108 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13280 62863
rect 13108 62759 13280 62817
rect 13108 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13280 62759
rect 13108 62655 13280 62713
rect 13108 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13280 62655
rect 13108 62551 13280 62609
rect 13108 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13280 62551
rect 13108 62447 13280 62505
rect 13108 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13280 62447
rect 13108 62343 13280 62401
rect 13108 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13280 62343
rect 13108 62239 13280 62297
rect 13108 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13280 62239
rect 13108 62135 13280 62193
rect 13108 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13280 62135
rect 13108 62031 13280 62089
rect 13108 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13280 62031
rect 13108 61927 13280 61985
rect 13108 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13280 61927
rect 13108 61823 13280 61881
rect 13108 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13280 61823
rect 13108 61719 13280 61777
rect 13108 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13280 61719
rect 13108 61615 13280 61673
rect 13108 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13280 61615
rect 13108 61511 13280 61569
rect 13108 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13280 61511
rect 13108 61407 13280 61465
rect 13108 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13280 61407
rect 13108 61303 13280 61361
rect 13108 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13280 61303
rect 13108 61199 13280 61257
rect 13108 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13280 61199
rect 13108 61095 13280 61153
rect 13108 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13280 61095
rect 13108 60991 13280 61049
rect 13108 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13280 60991
rect 13108 60887 13280 60945
rect 13108 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13280 60887
rect 13108 60783 13280 60841
rect 13108 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13280 60783
rect 13108 60679 13280 60737
rect 13108 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13280 60679
rect 13108 60575 13280 60633
rect 13108 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13280 60575
rect 13108 60471 13280 60529
rect 13108 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13280 60471
rect 13108 60367 13280 60425
rect 13108 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13280 60367
rect 13108 60263 13280 60321
rect 13108 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13280 60263
rect 13108 60159 13280 60217
rect 13108 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13280 60159
rect 13108 60055 13280 60113
rect 13108 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13280 60055
rect 13108 59951 13280 60009
rect 13108 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13280 59951
rect 13108 59847 13280 59905
rect 13108 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13280 59847
rect 13108 59743 13280 59801
rect 13108 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13280 59743
rect 13108 59639 13280 59697
rect 13108 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13280 59639
rect 13108 59535 13280 59593
rect 13108 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13280 59535
rect 13108 59431 13280 59489
rect 13108 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13280 59431
rect 13108 59327 13280 59385
rect 13108 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13280 59327
rect 13108 59223 13280 59281
rect 13108 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13280 59223
rect 13108 59119 13280 59177
rect 13108 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13280 59119
rect 13108 59015 13280 59073
rect 13108 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13280 59015
rect 13108 58911 13280 58969
rect 13108 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13280 58911
rect 13108 58807 13280 58865
rect 13108 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13280 58807
rect 13108 58703 13280 58761
rect 13108 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13280 58703
rect 13108 58599 13280 58657
rect 13108 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13280 58599
rect 13108 58495 13280 58553
rect 13108 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13280 58495
rect 13108 58391 13280 58449
rect 13108 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13280 58391
rect 13108 58287 13280 58345
rect 13108 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13280 58287
rect 13108 58183 13280 58241
rect 13108 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13280 58183
rect 13108 58079 13280 58137
rect 13108 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13280 58079
rect 13108 57975 13280 58033
rect 13108 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13280 57975
rect 13108 57871 13280 57929
rect 13108 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13280 57871
rect 13108 57767 13280 57825
rect 13108 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13280 57767
rect 13108 57663 13280 57721
rect 13108 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13280 57663
rect 13108 57559 13280 57617
rect 13108 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13280 57559
rect 13108 57455 13280 57513
rect 13108 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13280 57455
rect 13108 57351 13280 57409
rect 13108 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13280 57351
rect 13108 57247 13280 57305
rect 13108 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13280 57247
rect 13108 57143 13280 57201
rect 13108 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13280 57143
rect 13108 57039 13280 57097
rect 13108 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13280 57039
rect 13108 56935 13280 56993
rect 13108 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13280 56935
rect 13108 56831 13280 56889
rect 13108 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13280 56831
rect 13108 56727 13280 56785
rect 13108 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13280 56727
rect 13108 56623 13280 56681
rect 13108 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13280 56623
rect 13108 56519 13280 56577
rect 13108 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13280 56519
rect 13108 56415 13280 56473
rect 13108 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13280 56415
rect 13108 56311 13280 56369
rect 13108 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13280 56311
rect 13108 56207 13280 56265
rect 13108 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13280 56207
rect 13108 56103 13280 56161
rect 13108 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13280 56103
rect 13108 55999 13280 56057
rect 13108 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13280 55999
rect 13108 55895 13280 55953
rect 13108 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13280 55895
rect 13108 55791 13280 55849
rect 13108 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13280 55791
rect 13108 55687 13280 55745
rect 13108 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13280 55687
rect 13108 55583 13280 55641
rect 13108 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13280 55583
rect 13108 55479 13280 55537
rect 13108 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13280 55479
rect 13108 55375 13280 55433
rect 13108 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13280 55375
rect 13108 55271 13280 55329
rect 13108 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13280 55271
rect 13108 55167 13280 55225
rect 13108 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13280 55167
rect 13108 55063 13280 55121
rect 13108 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13280 55063
rect 13108 54959 13280 55017
rect 13108 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13280 54959
rect 13108 54855 13280 54913
rect 13108 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13280 54855
rect 13108 54751 13280 54809
rect 13108 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13280 54751
rect 13108 54647 13280 54705
rect 13108 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13280 54647
rect 13108 54543 13280 54601
rect 13108 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13280 54543
rect 13108 54439 13280 54497
rect 13108 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13280 54439
rect 13108 54335 13280 54393
rect 13108 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13280 54335
rect 13108 54231 13280 54289
rect 13108 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13280 54231
rect 13108 54127 13280 54185
rect 13108 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13280 54127
rect 13108 54023 13280 54081
rect 13108 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13280 54023
rect 13108 53919 13280 53977
rect 13108 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13280 53919
rect 13108 53815 13280 53873
rect 13108 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13280 53815
rect 13108 53711 13280 53769
rect 13108 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13280 53711
rect 13108 53607 13280 53665
rect 13108 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13280 53607
rect 13108 53503 13280 53561
rect 13108 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13280 53503
rect 13108 53399 13280 53457
rect 13108 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13280 53399
rect 13108 53295 13280 53353
rect 13108 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13280 53295
rect 13108 53191 13280 53249
rect 13108 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13280 53191
rect 13108 53087 13280 53145
rect 13108 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13280 53087
rect 13108 52983 13280 53041
rect 13108 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13280 52983
rect 13108 52879 13280 52937
rect 13108 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13280 52879
rect 13108 52775 13280 52833
rect 13108 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13280 52775
rect 13108 52671 13280 52729
rect 13108 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13280 52671
rect 13108 52567 13280 52625
rect 13108 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13280 52567
rect 13108 52463 13280 52521
rect 13108 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13280 52463
rect 13108 52359 13280 52417
rect 13108 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13280 52359
rect 13108 52255 13280 52313
rect 13108 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13280 52255
rect 13108 52151 13280 52209
rect 13108 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13280 52151
rect 13108 52047 13280 52105
rect 13108 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13280 52047
rect 13108 51943 13280 52001
rect 13108 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13280 51943
rect 13108 51839 13280 51897
rect 13108 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13280 51839
rect 13108 51735 13280 51793
rect 13108 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13280 51735
rect 13108 51631 13280 51689
rect 13108 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13280 51631
rect 13108 51527 13280 51585
rect 13108 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13280 51527
rect 13108 51423 13280 51481
rect 13108 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13280 51423
rect 13108 51319 13280 51377
rect 13108 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13280 51319
rect 13108 51215 13280 51273
rect 13108 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13280 51215
rect 13108 51111 13280 51169
rect 13108 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13280 51111
rect 13108 51007 13280 51065
rect 13108 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13280 51007
rect 13108 50903 13280 50961
rect 13108 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13280 50903
rect 13108 50799 13280 50857
rect 13108 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13280 50799
rect 13108 50695 13280 50753
rect 13108 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13280 50695
rect 13108 50591 13280 50649
rect 13108 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13280 50591
rect 13108 50487 13280 50545
rect 13108 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13280 50487
rect 13108 50383 13280 50441
rect 13108 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13280 50383
rect 13108 50279 13280 50337
rect 13108 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13280 50279
rect 13108 50175 13280 50233
rect 13108 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13280 50175
rect 13108 50071 13280 50129
rect 13108 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13280 50071
rect 13108 49967 13280 50025
rect 13108 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13280 49967
rect 13108 49863 13280 49921
rect 13108 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13280 49863
rect 13108 49759 13280 49817
rect 13108 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13280 49759
rect 13108 49655 13280 49713
rect 13108 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13280 49655
rect 13108 49551 13280 49609
rect 13108 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13280 49551
rect 13108 49447 13280 49505
rect 13108 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13280 49447
rect 13108 49343 13280 49401
rect 13108 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13280 49343
rect 13108 49239 13280 49297
rect 13108 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13280 49239
rect 13108 49135 13280 49193
rect 13108 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13280 49135
rect 13108 49031 13280 49089
rect 13108 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13280 49031
rect 13108 48927 13280 48985
rect 13108 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13280 48927
rect 13108 48823 13280 48881
rect 13108 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13280 48823
rect 13108 48719 13280 48777
rect 13108 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13280 48719
rect 13108 48615 13280 48673
rect 13108 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13280 48615
rect 13108 48511 13280 48569
rect 13108 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13280 48511
rect 13108 48407 13280 48465
rect 13108 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13280 48407
rect 13108 48303 13280 48361
rect 13108 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13280 48303
rect 13108 48199 13280 48257
rect 13108 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13280 48199
rect 13108 48095 13280 48153
rect 13108 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13280 48095
rect 13108 47991 13280 48049
rect 13108 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13280 47991
rect 13108 47887 13280 47945
rect 13108 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13280 47887
rect 13108 47783 13280 47841
rect 13108 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13280 47783
rect 13108 47679 13280 47737
rect 13108 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13280 47679
rect 13108 47575 13280 47633
rect 13108 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13280 47575
rect 13108 47471 13280 47529
rect 13108 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13280 47471
rect 13108 47367 13280 47425
rect 13108 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13280 47367
rect 13108 47263 13280 47321
rect 13108 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13280 47263
rect 13108 47159 13280 47217
rect 13108 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13280 47159
rect 13108 47055 13280 47113
rect 13108 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13280 47055
rect 13108 46951 13280 47009
rect 13108 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13280 46951
rect 13108 46847 13280 46905
rect 13108 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13280 46847
rect 13108 46743 13280 46801
rect 13108 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13280 46743
rect 13108 46639 13280 46697
rect 13108 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13280 46639
rect 13108 46535 13280 46593
rect 13108 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13280 46535
rect 13108 46431 13280 46489
rect 13108 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13280 46431
rect 13108 46327 13280 46385
rect 13108 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13280 46327
rect 13108 46223 13280 46281
rect 13108 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13280 46223
rect 13108 46119 13280 46177
rect 13108 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13280 46119
rect 13108 46015 13280 46073
rect 13108 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13280 46015
rect 13108 45911 13280 45969
rect 13108 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13280 45911
rect 13108 45807 13280 45865
rect 13108 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13280 45807
rect 13108 45703 13280 45761
rect 13108 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13280 45703
rect 13108 45599 13280 45657
rect 13108 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13280 45599
rect 13108 45495 13280 45553
rect 13108 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13280 45495
rect 13108 45391 13280 45449
rect 13108 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13280 45391
rect 13108 45287 13280 45345
rect 13108 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13280 45287
rect 13108 45183 13280 45241
rect 13108 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13280 45183
rect 13108 45079 13280 45137
rect 13108 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13280 45079
rect 13108 44902 13280 45033
rect 70813 69758 70824 69785
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70813 69700 71000 69758
rect 70813 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70813 69596 71000 69654
rect 70813 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70813 69492 71000 69550
rect 70813 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70813 69388 71000 69446
rect 70813 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70813 69284 71000 69342
rect 70813 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70813 69180 71000 69238
rect 70813 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70813 69076 71000 69134
rect 70813 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70813 68972 71000 69030
rect 70813 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70813 68868 71000 68926
rect 70813 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70813 68764 71000 68822
rect 70813 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70813 68660 71000 68718
rect 70813 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70813 68556 71000 68614
rect 70813 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70813 68452 71000 68510
rect 70813 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70813 68348 71000 68406
rect 70813 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70813 68244 71000 68302
rect 70813 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70813 68140 71000 68198
rect 70813 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70813 68036 71000 68094
rect 70813 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70813 67932 71000 67990
rect 70813 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70813 67828 71000 67886
rect 70813 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70813 67724 71000 67782
rect 70813 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70813 67620 71000 67678
rect 70813 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70813 67516 71000 67574
rect 70813 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70813 67412 71000 67470
rect 70813 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70813 67308 71000 67366
rect 70813 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70813 67204 71000 67262
rect 70813 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70813 67100 71000 67158
rect 70813 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70813 66996 71000 67054
rect 70813 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70813 66892 71000 66950
rect 70813 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70813 66788 71000 66846
rect 70813 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70813 66684 71000 66742
rect 70813 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70813 66580 71000 66638
rect 70813 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70813 66476 71000 66534
rect 70813 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70813 66372 71000 66430
rect 70813 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70813 66268 71000 66326
rect 70813 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70813 66164 71000 66222
rect 70813 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70813 66060 71000 66118
rect 70813 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70813 65956 71000 66014
rect 70813 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70813 65852 71000 65910
rect 70813 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70813 65748 71000 65806
rect 70813 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70813 65644 71000 65702
rect 70813 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70813 65540 71000 65598
rect 70813 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70813 65436 71000 65494
rect 70813 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70813 65332 71000 65390
rect 70813 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70813 65228 71000 65286
rect 70813 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70813 65124 71000 65182
rect 70813 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70813 65020 71000 65078
rect 70813 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70813 64916 71000 64974
rect 70813 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70813 64812 71000 64870
rect 70813 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70813 64708 71000 64766
rect 70813 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70813 64604 71000 64662
rect 70813 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70813 64500 71000 64558
rect 70813 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70813 64396 71000 64454
rect 70813 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70813 64292 71000 64350
rect 70813 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70813 64188 71000 64246
rect 70813 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70813 64084 71000 64142
rect 70813 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70813 63980 71000 64038
rect 70813 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70813 63876 71000 63934
rect 70813 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70813 63772 71000 63830
rect 70813 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70813 63668 71000 63726
rect 70813 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70813 63564 71000 63622
rect 70813 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70813 63460 71000 63518
rect 70813 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70813 63356 71000 63414
rect 70813 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70813 63252 71000 63310
rect 70813 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70813 63148 71000 63206
rect 70813 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70813 63044 71000 63102
rect 70813 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70813 62940 71000 62998
rect 70813 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70813 62836 71000 62894
rect 70813 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70813 62732 71000 62790
rect 70813 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70813 62628 71000 62686
rect 70813 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70813 62524 71000 62582
rect 70813 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70813 62420 71000 62478
rect 70813 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70813 62316 71000 62374
rect 70813 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70813 62212 71000 62270
rect 70813 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70813 62108 71000 62166
rect 70813 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70813 62004 71000 62062
rect 70813 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70813 61900 71000 61958
rect 70813 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70813 61796 71000 61854
rect 70813 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70813 61692 71000 61750
rect 70813 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70813 61588 71000 61646
rect 70813 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70813 61484 71000 61542
rect 70813 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70813 61380 71000 61438
rect 70813 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70813 61276 71000 61334
rect 70813 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70813 61172 71000 61230
rect 70813 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70813 61068 71000 61126
rect 70813 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70813 60964 71000 61022
rect 70813 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70813 60860 71000 60918
rect 70813 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70813 60756 71000 60814
rect 70813 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70813 60652 71000 60710
rect 70813 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70813 60548 71000 60606
rect 70813 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70813 60444 71000 60502
rect 70813 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70813 60340 71000 60398
rect 70813 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70813 60236 71000 60294
rect 70813 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70813 60132 71000 60190
rect 70813 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70813 60028 71000 60086
rect 70813 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70813 59924 71000 59982
rect 70813 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70813 59820 71000 59878
rect 70813 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70813 59716 71000 59774
rect 70813 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70813 59612 71000 59670
rect 70813 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70813 59508 71000 59566
rect 70813 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70813 59404 71000 59462
rect 70813 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70813 59300 71000 59358
rect 70813 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70813 59196 71000 59254
rect 70813 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70813 59092 71000 59150
rect 70813 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70813 58988 71000 59046
rect 70813 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70813 58884 71000 58942
rect 70813 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70813 58780 71000 58838
rect 70813 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70813 58676 71000 58734
rect 70813 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70813 58572 71000 58630
rect 70813 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70813 58468 71000 58526
rect 70813 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70813 58364 71000 58422
rect 70813 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70813 58260 71000 58318
rect 70813 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70813 58156 71000 58214
rect 70813 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70813 58052 71000 58110
rect 70813 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70813 57948 71000 58006
rect 70813 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70813 57844 71000 57902
rect 70813 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70813 57740 71000 57798
rect 70813 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70813 57636 71000 57694
rect 70813 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70813 57532 71000 57590
rect 70813 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70813 57428 71000 57486
rect 70813 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70813 57324 71000 57382
rect 70813 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70813 57220 71000 57278
rect 70813 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70813 57116 71000 57174
rect 70813 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70813 57012 71000 57070
rect 70813 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70813 56908 71000 56966
rect 70813 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70813 56804 71000 56862
rect 70813 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70813 56700 71000 56758
rect 70813 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70813 56596 71000 56654
rect 70813 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70813 56492 71000 56550
rect 70813 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70813 56388 71000 56446
rect 70813 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70813 56284 71000 56342
rect 70813 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70813 56180 71000 56238
rect 70813 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70813 56076 71000 56134
rect 70813 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70813 55972 71000 56030
rect 70813 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70813 55868 71000 55926
rect 70813 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70813 55764 71000 55822
rect 70813 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70813 55660 71000 55718
rect 70813 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70813 55556 71000 55614
rect 70813 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70813 55452 71000 55510
rect 70813 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70813 55348 71000 55406
rect 70813 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70813 55244 71000 55302
rect 70813 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70813 55140 71000 55198
rect 70813 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70813 55036 71000 55094
rect 70813 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70813 54932 71000 54990
rect 70813 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70813 54828 71000 54886
rect 70813 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70813 54724 71000 54782
rect 70813 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70813 54620 71000 54678
rect 70813 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70813 54516 71000 54574
rect 70813 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70813 54412 71000 54470
rect 70813 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70813 54308 71000 54366
rect 70813 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70813 54204 71000 54262
rect 70813 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70813 54100 71000 54158
rect 70813 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70813 53996 71000 54054
rect 70813 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70813 53892 71000 53950
rect 70813 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70813 53788 71000 53846
rect 70813 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70813 53684 71000 53742
rect 70813 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70813 53580 71000 53638
rect 70813 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70813 53476 71000 53534
rect 70813 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70813 53372 71000 53430
rect 70813 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70813 53268 71000 53326
rect 70813 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70813 53164 71000 53222
rect 70813 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70813 53060 71000 53118
rect 70813 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70813 52956 71000 53014
rect 70813 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70813 52852 71000 52910
rect 70813 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70813 52748 71000 52806
rect 70813 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70813 52644 71000 52702
rect 70813 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70813 52540 71000 52598
rect 70813 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70813 52436 71000 52494
rect 70813 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70813 52332 71000 52390
rect 70813 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70813 52228 71000 52286
rect 70813 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70813 52124 71000 52182
rect 70813 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70813 52020 71000 52078
rect 70813 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70813 51916 71000 51974
rect 70813 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70813 51812 71000 51870
rect 70813 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70813 51708 71000 51766
rect 70813 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70813 51604 71000 51662
rect 70813 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70813 51500 71000 51558
rect 70813 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70813 51396 71000 51454
rect 70813 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70813 51292 71000 51350
rect 70813 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70813 51188 71000 51246
rect 70813 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70813 51084 71000 51142
rect 70813 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70813 50980 71000 51038
rect 70813 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70813 50876 71000 50934
rect 70813 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70813 50772 71000 50830
rect 70813 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70813 50668 71000 50726
rect 70813 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70813 50564 71000 50622
rect 70813 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70813 50460 71000 50518
rect 70813 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70813 50356 71000 50414
rect 70813 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70813 50252 71000 50310
rect 70813 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70813 50148 71000 50206
rect 70813 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70813 50044 71000 50102
rect 70813 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70813 49940 71000 49998
rect 70813 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70813 49836 71000 49894
rect 70813 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70813 49732 71000 49790
rect 70813 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70813 49628 71000 49686
rect 70813 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70813 49524 71000 49582
rect 70813 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70813 49420 71000 49478
rect 70813 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70813 49316 71000 49374
rect 70813 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70813 49212 71000 49270
rect 70813 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70813 49108 71000 49166
rect 70813 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70813 49004 71000 49062
rect 70813 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70813 48900 71000 48958
rect 70813 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70813 48796 71000 48854
rect 70813 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70813 48692 71000 48750
rect 70813 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70813 48588 71000 48646
rect 70813 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70813 48484 71000 48542
rect 70813 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70813 48380 71000 48438
rect 70813 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70813 48276 71000 48334
rect 70813 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70813 48172 71000 48230
rect 70813 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70813 48068 71000 48126
rect 70813 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70813 47964 71000 48022
rect 70813 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70813 47860 71000 47918
rect 70813 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70813 47756 71000 47814
rect 70813 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70813 47652 71000 47710
rect 70813 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70813 47548 71000 47606
rect 70813 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70813 47444 71000 47502
rect 70813 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70813 47340 71000 47398
rect 70813 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70813 47236 71000 47294
rect 70813 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70813 47132 71000 47190
rect 70813 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70813 47028 71000 47086
rect 70813 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70813 46924 71000 46982
rect 70813 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70813 46820 71000 46878
rect 70813 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70813 46716 71000 46774
rect 70813 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70813 46612 71000 46670
rect 70813 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70813 46508 71000 46566
rect 70813 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70813 46404 71000 46462
rect 70813 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70813 46300 71000 46358
rect 70813 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70813 46196 71000 46254
rect 70813 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70813 46092 71000 46150
rect 70813 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70813 45988 71000 46046
rect 70813 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70813 45884 71000 45942
rect 70813 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70813 45780 71000 45838
rect 70813 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70813 45676 71000 45734
rect 70813 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70813 45572 71000 45630
rect 70813 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70813 45468 71000 45526
rect 70813 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70813 45364 71000 45422
rect 70813 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70813 45260 71000 45318
rect 70813 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70813 45156 71000 45214
rect 70813 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70813 45052 71000 45110
rect 70813 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70813 44948 71000 45006
tri 13280 44902 13298 44920 sw
rect 70813 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13108 44848 13298 44902
tri 13108 44844 13112 44848 ne
rect 13112 44844 13298 44848
tri 13298 44844 13356 44902 sw
rect 70813 44844 71000 44902
tri 13112 44824 13132 44844 ne
rect 13132 44824 13356 44844
tri 13356 44824 13376 44844 sw
tri 13132 44778 13178 44824 ne
rect 13178 44778 13254 44824
rect 13300 44798 13376 44824
tri 13376 44798 13402 44824 sw
rect 70813 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 13300 44778 13402 44798
tri 13402 44778 13422 44798 sw
tri 13178 44740 13216 44778 ne
rect 13216 44740 13422 44778
tri 13422 44740 13460 44778 sw
rect 70813 44740 71000 44798
tri 13216 44694 13262 44740 ne
rect 13262 44694 13460 44740
tri 13460 44694 13506 44740 sw
rect 70813 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
tri 13262 44692 13264 44694 ne
rect 13264 44692 13506 44694
tri 13506 44692 13508 44694 sw
tri 13264 44646 13310 44692 ne
rect 13310 44646 13386 44692
rect 13432 44646 13508 44692
tri 13310 44636 13320 44646 ne
rect 13320 44636 13508 44646
tri 13508 44636 13564 44692 sw
rect 70813 44636 71000 44694
tri 13320 44590 13366 44636 ne
rect 13366 44590 13564 44636
tri 13564 44590 13610 44636 sw
rect 70813 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13366 44560 13396 44590 ne
rect 13396 44560 13610 44590
tri 13610 44560 13640 44590 sw
tri 13396 44514 13442 44560 ne
rect 13442 44514 13518 44560
rect 13564 44532 13640 44560
tri 13640 44532 13668 44560 sw
rect 70813 44532 71000 44590
rect 13564 44514 13668 44532
tri 13668 44514 13686 44532 sw
tri 13442 44486 13470 44514 ne
rect 13470 44486 13686 44514
tri 13686 44486 13714 44514 sw
rect 70813 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
tri 13470 44428 13528 44486 ne
rect 13528 44428 13714 44486
tri 13714 44428 13772 44486 sw
rect 70813 44428 71000 44486
tri 13528 44382 13574 44428 ne
rect 13574 44382 13650 44428
rect 13696 44382 13772 44428
tri 13772 44382 13818 44428 sw
rect 70813 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
tri 13574 44324 13632 44382 ne
rect 13632 44324 13818 44382
tri 13818 44324 13876 44382 sw
rect 70813 44324 71000 44382
tri 13632 44296 13660 44324 ne
rect 13660 44296 13876 44324
tri 13876 44296 13904 44324 sw
tri 13660 44250 13706 44296 ne
rect 13706 44250 13782 44296
rect 13828 44278 13904 44296
tri 13904 44278 13922 44296 sw
rect 70813 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 13828 44250 13922 44278
tri 13706 44220 13736 44250 ne
rect 13736 44220 13922 44250
tri 13922 44220 13980 44278 sw
rect 70813 44220 71000 44278
tri 13736 44174 13782 44220 ne
rect 13782 44174 13980 44220
tri 13980 44174 14026 44220 sw
rect 70813 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
tri 13782 44164 13792 44174 ne
rect 13792 44164 14026 44174
tri 14026 44164 14036 44174 sw
tri 13792 44118 13838 44164 ne
rect 13838 44118 13914 44164
rect 13960 44118 14036 44164
tri 14036 44118 14082 44164 sw
tri 13838 44116 13840 44118 ne
rect 13840 44116 14082 44118
tri 14082 44116 14084 44118 sw
rect 70813 44116 71000 44174
tri 13840 44070 13886 44116 ne
rect 13886 44070 14084 44116
tri 14084 44070 14130 44116 sw
rect 70813 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
tri 13886 44032 13924 44070 ne
rect 13924 44032 14130 44070
tri 13924 43986 13970 44032 ne
rect 13970 43986 14046 44032
rect 14092 44012 14130 44032
tri 14130 44012 14188 44070 sw
rect 70813 44012 71000 44070
rect 14092 43986 14188 44012
tri 13970 43966 13990 43986 ne
rect 13990 43966 14188 43986
tri 14188 43966 14234 44012 sw
rect 70813 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13990 43908 14048 43966 ne
rect 14048 43908 14234 43966
tri 14234 43908 14292 43966 sw
rect 70813 43908 71000 43966
tri 14048 43900 14056 43908 ne
rect 14056 43900 14292 43908
tri 14292 43900 14300 43908 sw
tri 14056 43854 14102 43900 ne
rect 14102 43854 14178 43900
rect 14224 43862 14300 43900
tri 14300 43862 14338 43900 sw
rect 70813 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 14224 43854 14338 43862
tri 14102 43852 14104 43854 ne
rect 14104 43852 14338 43854
tri 14104 43804 14152 43852 ne
rect 14152 43804 14338 43852
tri 14338 43804 14396 43862 sw
rect 70813 43804 71000 43862
tri 14152 43768 14188 43804 ne
rect 14188 43768 14396 43804
tri 14396 43768 14432 43804 sw
tri 14188 43722 14234 43768 ne
rect 14234 43722 14310 43768
rect 14356 43758 14432 43768
tri 14432 43758 14442 43768 sw
rect 70813 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43722 14442 43758
tri 14442 43722 14478 43758 sw
tri 14234 43700 14256 43722 ne
rect 14256 43700 14478 43722
tri 14478 43700 14500 43722 sw
rect 70813 43700 71000 43758
tri 14256 43654 14302 43700 ne
rect 14302 43654 14500 43700
tri 14500 43654 14546 43700 sw
rect 70813 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
tri 14302 43636 14320 43654 ne
rect 14320 43636 14546 43654
tri 14546 43636 14564 43654 sw
tri 14320 43590 14366 43636 ne
rect 14366 43590 14442 43636
rect 14488 43596 14564 43636
tri 14564 43596 14604 43636 sw
rect 70813 43596 71000 43654
rect 14488 43590 14604 43596
tri 14366 43550 14406 43590 ne
rect 14406 43550 14604 43590
tri 14604 43550 14650 43596 sw
rect 70813 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
tri 14406 43504 14452 43550 ne
rect 14452 43504 14650 43550
tri 14650 43504 14696 43550 sw
tri 14452 43458 14498 43504 ne
rect 14498 43458 14574 43504
rect 14620 43492 14696 43504
tri 14696 43492 14708 43504 sw
rect 70813 43492 71000 43550
rect 14620 43458 14708 43492
tri 14708 43458 14742 43492 sw
tri 14498 43446 14510 43458 ne
rect 14510 43446 14742 43458
tri 14742 43446 14754 43458 sw
rect 70813 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14510 43388 14568 43446 ne
rect 14568 43388 14754 43446
tri 14754 43388 14812 43446 sw
rect 70813 43388 71000 43446
tri 14568 43372 14584 43388 ne
rect 14584 43372 14812 43388
tri 14584 43326 14630 43372 ne
rect 14630 43326 14706 43372
rect 14752 43342 14812 43372
tri 14812 43342 14858 43388 sw
rect 70813 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 14752 43326 14858 43342
tri 14630 43284 14672 43326 ne
rect 14672 43284 14858 43326
tri 14858 43284 14916 43342 sw
rect 70813 43284 71000 43342
tri 14672 43240 14716 43284 ne
rect 14716 43240 14916 43284
tri 14916 43240 14960 43284 sw
tri 14716 43194 14762 43240 ne
rect 14762 43194 14838 43240
rect 14884 43238 14960 43240
tri 14960 43238 14962 43240 sw
rect 70813 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43194 14962 43238
tri 14762 43180 14776 43194 ne
rect 14776 43180 14962 43194
tri 14962 43180 15020 43238 sw
rect 70813 43180 71000 43238
tri 14776 43134 14822 43180 ne
rect 14822 43134 15020 43180
tri 15020 43134 15066 43180 sw
rect 70813 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14822 43108 14848 43134 ne
rect 14848 43108 15066 43134
tri 15066 43108 15092 43134 sw
tri 14848 43062 14894 43108 ne
rect 14894 43062 14970 43108
rect 15016 43076 15092 43108
tri 15092 43076 15124 43108 sw
rect 70813 43076 71000 43134
rect 15016 43062 15124 43076
tri 15124 43062 15138 43076 sw
tri 14894 43030 14926 43062 ne
rect 14926 43030 15138 43062
tri 15138 43030 15170 43062 sw
rect 70813 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14926 42976 14980 43030 ne
rect 14980 42976 15170 43030
tri 14980 42930 15026 42976 ne
rect 15026 42930 15102 42976
rect 15148 42972 15170 42976
tri 15170 42972 15228 43030 sw
rect 70813 42972 71000 43030
rect 15148 42930 15228 42972
tri 15026 42926 15030 42930 ne
rect 15030 42926 15228 42930
tri 15228 42926 15274 42972 sw
rect 70813 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15030 42868 15088 42926 ne
rect 15088 42868 15274 42926
tri 15274 42868 15332 42926 sw
rect 70813 42868 71000 42926
tri 15088 42844 15112 42868 ne
rect 15112 42844 15332 42868
tri 15332 42844 15356 42868 sw
tri 15112 42798 15158 42844 ne
rect 15158 42798 15234 42844
rect 15280 42822 15356 42844
tri 15356 42822 15378 42844 sw
rect 70813 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 15280 42798 15378 42822
tri 15158 42764 15192 42798 ne
rect 15192 42764 15378 42798
tri 15378 42764 15436 42822 sw
rect 70813 42764 71000 42822
tri 15192 42718 15238 42764 ne
rect 15238 42718 15436 42764
tri 15436 42718 15482 42764 sw
rect 70813 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
tri 15238 42712 15244 42718 ne
rect 15244 42712 15482 42718
tri 15482 42712 15488 42718 sw
tri 15244 42666 15290 42712 ne
rect 15290 42666 15366 42712
rect 15412 42666 15488 42712
tri 15488 42666 15534 42712 sw
tri 15290 42660 15296 42666 ne
rect 15296 42660 15534 42666
tri 15534 42660 15540 42666 sw
rect 70813 42660 71000 42718
tri 15296 42614 15342 42660 ne
rect 15342 42614 15540 42660
tri 15540 42614 15586 42660 sw
rect 70813 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15342 42580 15376 42614 ne
rect 15376 42580 15586 42614
tri 15376 42534 15422 42580 ne
rect 15422 42534 15498 42580
rect 15544 42556 15586 42580
tri 15586 42556 15644 42614 sw
rect 70813 42556 71000 42614
rect 15544 42534 15644 42556
tri 15422 42510 15446 42534 ne
rect 15446 42510 15644 42534
tri 15644 42510 15690 42556 sw
rect 70813 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
tri 15446 42452 15504 42510 ne
rect 15504 42452 15690 42510
tri 15690 42452 15748 42510 sw
rect 70813 42452 71000 42510
tri 15504 42448 15508 42452 ne
rect 15508 42448 15748 42452
tri 15748 42448 15752 42452 sw
tri 15508 42402 15554 42448 ne
rect 15554 42402 15630 42448
rect 15676 42406 15752 42448
tri 15752 42406 15794 42448 sw
rect 70813 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 15676 42402 15794 42406
tri 15554 42388 15568 42402 ne
rect 15568 42388 15794 42402
tri 15568 42348 15608 42388 ne
rect 15608 42348 15794 42388
tri 15794 42348 15852 42406 sw
rect 70813 42348 71000 42406
tri 15608 42316 15640 42348 ne
rect 15640 42316 15852 42348
tri 15852 42316 15884 42348 sw
tri 15640 42270 15686 42316 ne
rect 15686 42270 15762 42316
rect 15808 42302 15884 42316
tri 15884 42302 15898 42316 sw
rect 70813 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42270 15898 42302
tri 15898 42270 15930 42302 sw
tri 15686 42244 15712 42270 ne
rect 15712 42244 15930 42270
tri 15930 42244 15956 42270 sw
rect 70813 42244 71000 42302
tri 15712 42198 15758 42244 ne
rect 15758 42198 15956 42244
tri 15956 42198 16002 42244 sw
rect 70813 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
tri 15758 42184 15772 42198 ne
rect 15772 42184 16002 42198
tri 16002 42184 16016 42198 sw
tri 15772 42138 15818 42184 ne
rect 15818 42138 15894 42184
rect 15940 42140 16016 42184
tri 16016 42140 16060 42184 sw
rect 70813 42140 71000 42198
rect 15940 42138 16060 42140
tri 15818 42094 15862 42138 ne
rect 15862 42094 16060 42138
tri 16060 42094 16106 42140 sw
rect 70813 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15862 42052 15904 42094 ne
rect 15904 42052 16106 42094
tri 16106 42052 16148 42094 sw
tri 15904 42006 15950 42052 ne
rect 15950 42006 16026 42052
rect 16072 42036 16148 42052
tri 16148 42036 16164 42052 sw
rect 70813 42036 71000 42094
rect 16072 42006 16164 42036
tri 16164 42006 16194 42036 sw
tri 15950 41990 15966 42006 ne
rect 15966 41990 16194 42006
tri 16194 41990 16210 42006 sw
rect 70813 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15966 41932 16024 41990 ne
rect 16024 41932 16210 41990
tri 16210 41932 16268 41990 sw
rect 70813 41932 71000 41990
tri 16024 41920 16036 41932 ne
rect 16036 41920 16268 41932
tri 16036 41874 16082 41920 ne
rect 16082 41874 16158 41920
rect 16204 41886 16268 41920
tri 16268 41886 16314 41932 sw
rect 70813 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 16204 41874 16314 41886
tri 16082 41828 16128 41874 ne
rect 16128 41828 16314 41874
tri 16314 41828 16372 41886 sw
rect 70813 41828 71000 41886
tri 16128 41788 16168 41828 ne
rect 16168 41788 16372 41828
tri 16372 41788 16412 41828 sw
tri 16168 41742 16214 41788 ne
rect 16214 41742 16290 41788
rect 16336 41782 16412 41788
tri 16412 41782 16418 41788 sw
rect 70813 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41742 16418 41782
tri 16214 41724 16232 41742 ne
rect 16232 41724 16418 41742
tri 16418 41724 16476 41782 sw
rect 70813 41724 71000 41782
tri 16232 41678 16278 41724 ne
rect 16278 41678 16476 41724
tri 16476 41678 16522 41724 sw
rect 70813 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
tri 16278 41656 16300 41678 ne
rect 16300 41656 16522 41678
tri 16522 41656 16544 41678 sw
tri 16300 41610 16346 41656 ne
rect 16346 41610 16422 41656
rect 16468 41620 16544 41656
tri 16544 41620 16580 41656 sw
rect 70813 41620 71000 41678
rect 16468 41610 16580 41620
tri 16580 41610 16590 41620 sw
tri 16346 41574 16382 41610 ne
rect 16382 41574 16590 41610
tri 16590 41574 16626 41610 sw
rect 70813 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16382 41524 16432 41574 ne
rect 16432 41524 16626 41574
tri 16432 41478 16478 41524 ne
rect 16478 41478 16554 41524
rect 16600 41516 16626 41524
tri 16626 41516 16684 41574 sw
rect 70813 41516 71000 41574
rect 16600 41478 16684 41516
tri 16478 41470 16486 41478 ne
rect 16486 41470 16684 41478
tri 16684 41470 16730 41516 sw
rect 70813 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
tri 16486 41412 16544 41470 ne
rect 16544 41412 16730 41470
tri 16730 41412 16788 41470 sw
rect 70813 41412 71000 41470
tri 16544 41392 16564 41412 ne
rect 16564 41392 16788 41412
tri 16788 41392 16808 41412 sw
tri 16564 41346 16610 41392 ne
rect 16610 41346 16686 41392
rect 16732 41366 16808 41392
tri 16808 41366 16834 41392 sw
rect 70813 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 16732 41346 16834 41366
tri 16610 41308 16648 41346 ne
rect 16648 41308 16834 41346
tri 16834 41308 16892 41366 sw
rect 70813 41308 71000 41366
tri 16648 41262 16694 41308 ne
rect 16694 41262 16892 41308
tri 16892 41262 16938 41308 sw
rect 70813 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
tri 16694 41260 16696 41262 ne
rect 16696 41260 16938 41262
tri 16938 41260 16940 41262 sw
tri 16696 41214 16742 41260 ne
rect 16742 41214 16818 41260
rect 16864 41214 16940 41260
tri 16940 41214 16986 41260 sw
tri 16742 41204 16752 41214 ne
rect 16752 41204 16986 41214
tri 16986 41204 16996 41214 sw
rect 70813 41204 71000 41262
tri 16752 41158 16798 41204 ne
rect 16798 41158 16996 41204
tri 16996 41158 17042 41204 sw
rect 70813 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
tri 16798 41128 16828 41158 ne
rect 16828 41128 17042 41158
tri 16828 41082 16874 41128 ne
rect 16874 41082 16950 41128
rect 16996 41100 17042 41128
tri 17042 41100 17100 41158 sw
rect 70813 41100 71000 41158
rect 16996 41082 17100 41100
tri 16874 41054 16902 41082 ne
rect 16902 41054 17100 41082
tri 17100 41054 17146 41100 sw
rect 70813 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
tri 16902 40996 16960 41054 ne
rect 16960 40996 17146 41054
tri 17146 40996 17204 41054 sw
rect 70813 40996 71000 41054
tri 16960 40950 17006 40996 ne
rect 17006 40950 17082 40996
rect 17128 40950 17204 40996
tri 17204 40950 17250 40996 sw
rect 70813 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
tri 17006 40924 17032 40950 ne
rect 17032 40924 17250 40950
tri 17032 40892 17064 40924 ne
rect 17064 40892 17250 40924
tri 17250 40892 17308 40950 sw
rect 70813 40892 71000 40950
tri 17064 40864 17092 40892 ne
rect 17092 40864 17308 40892
tri 17308 40864 17336 40892 sw
tri 17092 40818 17138 40864 ne
rect 17138 40818 17214 40864
rect 17260 40846 17336 40864
tri 17336 40846 17354 40864 sw
rect 70813 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40818 17354 40846
tri 17354 40818 17382 40846 sw
tri 17138 40788 17168 40818 ne
rect 17168 40788 17382 40818
tri 17382 40788 17412 40818 sw
rect 70813 40788 71000 40846
tri 17168 40742 17214 40788 ne
rect 17214 40742 17412 40788
tri 17412 40742 17458 40788 sw
rect 70813 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
tri 17214 40732 17224 40742 ne
rect 17224 40732 17458 40742
tri 17458 40732 17468 40742 sw
tri 17224 40686 17270 40732 ne
rect 17270 40686 17346 40732
rect 17392 40686 17468 40732
tri 17270 40684 17272 40686 ne
rect 17272 40684 17468 40686
tri 17468 40684 17516 40732 sw
rect 70813 40684 71000 40742
tri 17272 40638 17318 40684 ne
rect 17318 40638 17516 40684
tri 17516 40638 17562 40684 sw
rect 70813 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17318 40600 17356 40638 ne
rect 17356 40600 17562 40638
tri 17562 40600 17600 40638 sw
tri 17356 40554 17402 40600 ne
rect 17402 40554 17478 40600
rect 17524 40580 17600 40600
tri 17600 40580 17620 40600 sw
rect 70813 40580 71000 40638
rect 17524 40554 17620 40580
tri 17620 40554 17646 40580 sw
tri 17402 40534 17422 40554 ne
rect 17422 40534 17646 40554
tri 17646 40534 17666 40554 sw
rect 70813 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17422 40476 17480 40534 ne
rect 17480 40476 17666 40534
tri 17666 40476 17724 40534 sw
rect 70813 40476 71000 40534
tri 17480 40468 17488 40476 ne
rect 17488 40468 17724 40476
tri 17488 40422 17534 40468 ne
rect 17534 40422 17610 40468
rect 17656 40430 17724 40468
tri 17724 40430 17770 40476 sw
rect 70813 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 17656 40422 17770 40430
tri 17534 40372 17584 40422 ne
rect 17584 40372 17770 40422
tri 17770 40372 17828 40430 sw
rect 70813 40372 71000 40430
tri 17584 40336 17620 40372 ne
rect 17620 40336 17828 40372
tri 17828 40336 17864 40372 sw
tri 17620 40290 17666 40336 ne
rect 17666 40290 17742 40336
rect 17788 40326 17864 40336
tri 17864 40326 17874 40336 sw
rect 70813 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17788 40290 17874 40326
tri 17666 40268 17688 40290 ne
rect 17688 40268 17874 40290
tri 17874 40268 17932 40326 sw
rect 70813 40268 71000 40326
tri 17688 40222 17734 40268 ne
rect 17734 40222 17932 40268
tri 17932 40222 17978 40268 sw
rect 70813 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
tri 17734 40204 17752 40222 ne
rect 17752 40204 17978 40222
tri 17978 40204 17996 40222 sw
tri 17752 40158 17798 40204 ne
rect 17798 40158 17874 40204
rect 17920 40164 17996 40204
tri 17996 40164 18036 40204 sw
rect 70813 40164 71000 40222
rect 17920 40158 18036 40164
tri 18036 40158 18042 40164 sw
tri 17798 40118 17838 40158 ne
rect 17838 40118 18042 40158
tri 18042 40118 18082 40158 sw
rect 70813 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17838 40072 17884 40118 ne
rect 17884 40072 18082 40118
tri 17884 40026 17930 40072 ne
rect 17930 40026 18006 40072
rect 18052 40060 18082 40072
tri 18082 40060 18140 40118 sw
rect 70813 40060 71000 40118
rect 18052 40026 18140 40060
tri 17930 40014 17942 40026 ne
rect 17942 40014 18140 40026
tri 18140 40014 18186 40060 sw
rect 70813 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
tri 17942 39956 18000 40014 ne
rect 18000 39956 18186 40014
tri 18186 39956 18244 40014 sw
rect 70813 39956 71000 40014
tri 18000 39940 18016 39956 ne
rect 18016 39940 18244 39956
tri 18244 39940 18260 39956 sw
tri 18016 39894 18062 39940 ne
rect 18062 39894 18138 39940
rect 18184 39910 18260 39940
tri 18260 39910 18290 39940 sw
rect 70813 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 18184 39894 18290 39910
tri 18062 39852 18104 39894 ne
rect 18104 39852 18290 39894
tri 18290 39852 18348 39910 sw
rect 70813 39852 71000 39910
tri 18104 39808 18148 39852 ne
rect 18148 39808 18348 39852
tri 18348 39808 18392 39852 sw
tri 18148 39762 18194 39808 ne
rect 18194 39762 18270 39808
rect 18316 39806 18392 39808
tri 18392 39806 18394 39808 sw
rect 70813 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39762 18394 39806
tri 18394 39762 18438 39806 sw
tri 18194 39748 18208 39762 ne
rect 18208 39748 18438 39762
tri 18438 39748 18452 39762 sw
rect 70813 39748 71000 39806
tri 18208 39702 18254 39748 ne
rect 18254 39702 18452 39748
tri 18452 39702 18498 39748 sw
rect 70813 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
tri 18254 39676 18280 39702 ne
rect 18280 39676 18498 39702
tri 18280 39630 18326 39676 ne
rect 18326 39630 18402 39676
rect 18448 39644 18498 39676
tri 18498 39644 18556 39702 sw
rect 70813 39644 71000 39702
rect 18448 39630 18556 39644
tri 18326 39598 18358 39630 ne
rect 18358 39598 18556 39630
tri 18556 39598 18602 39644 sw
rect 70813 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18358 39544 18412 39598 ne
rect 18412 39544 18602 39598
tri 18602 39544 18656 39598 sw
tri 18412 39498 18458 39544 ne
rect 18458 39498 18534 39544
rect 18580 39540 18656 39544
tri 18656 39540 18660 39544 sw
rect 70813 39540 71000 39598
rect 18580 39498 18660 39540
tri 18660 39498 18702 39540 sw
tri 18458 39494 18462 39498 ne
rect 18462 39494 18702 39498
tri 18702 39494 18706 39498 sw
rect 70813 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18462 39460 18496 39494 ne
rect 18496 39460 18706 39494
tri 18496 39436 18520 39460 ne
rect 18520 39436 18706 39460
tri 18706 39436 18764 39494 sw
rect 70813 39436 71000 39494
tri 18520 39412 18544 39436 ne
rect 18544 39412 18764 39436
tri 18764 39412 18788 39436 sw
tri 18544 39366 18590 39412 ne
rect 18590 39366 18666 39412
rect 18712 39390 18788 39412
tri 18788 39390 18810 39412 sw
rect 70813 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 18712 39366 18810 39390
tri 18810 39366 18834 39390 sw
tri 18590 39332 18624 39366 ne
rect 18624 39332 18834 39366
tri 18834 39332 18868 39366 sw
rect 70813 39332 71000 39390
tri 18624 39286 18670 39332 ne
rect 18670 39286 18868 39332
tri 18868 39286 18914 39332 sw
rect 70813 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
tri 18670 39280 18676 39286 ne
rect 18676 39280 18914 39286
tri 18914 39280 18920 39286 sw
tri 18676 39234 18722 39280 ne
rect 18722 39234 18798 39280
rect 18844 39234 18920 39280
tri 18722 39228 18728 39234 ne
rect 18728 39228 18920 39234
tri 18920 39228 18972 39280 sw
rect 70813 39228 71000 39286
tri 18728 39182 18774 39228 ne
rect 18774 39182 18972 39228
tri 18972 39182 19018 39228 sw
rect 70813 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
tri 18774 39148 18808 39182 ne
rect 18808 39148 19018 39182
tri 19018 39148 19052 39182 sw
tri 18808 39102 18854 39148 ne
rect 18854 39102 18930 39148
rect 18976 39124 19052 39148
tri 19052 39124 19076 39148 sw
rect 70813 39124 71000 39182
rect 18976 39102 19076 39124
tri 19076 39102 19098 39124 sw
tri 18854 39078 18878 39102 ne
rect 18878 39078 19098 39102
tri 19098 39078 19122 39102 sw
rect 70813 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18878 39020 18936 39078 ne
rect 18936 39020 19122 39078
tri 19122 39020 19180 39078 sw
rect 70813 39020 71000 39078
tri 18936 39016 18940 39020 ne
rect 18940 39016 19180 39020
tri 18940 38970 18986 39016 ne
rect 18986 38970 19062 39016
rect 19108 38974 19180 39016
tri 19180 38974 19226 39020 sw
rect 70813 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 19108 38970 19226 38974
tri 18986 38916 19040 38970 ne
rect 19040 38916 19226 38970
tri 19226 38916 19284 38974 sw
rect 70813 38916 71000 38974
tri 19040 38884 19072 38916 ne
rect 19072 38884 19284 38916
tri 19284 38884 19316 38916 sw
tri 19072 38838 19118 38884 ne
rect 19118 38838 19194 38884
rect 19240 38870 19316 38884
tri 19316 38870 19330 38884 sw
rect 70813 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38838 19330 38870
tri 19118 38812 19144 38838 ne
rect 19144 38812 19330 38838
tri 19330 38812 19388 38870 sw
rect 70813 38812 71000 38870
tri 19144 38766 19190 38812 ne
rect 19190 38766 19388 38812
tri 19388 38766 19434 38812 sw
rect 70813 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19190 38752 19204 38766 ne
rect 19204 38752 19434 38766
tri 19434 38752 19448 38766 sw
tri 19204 38706 19250 38752 ne
rect 19250 38706 19326 38752
rect 19372 38708 19448 38752
tri 19448 38708 19492 38752 sw
rect 70813 38708 71000 38766
rect 19372 38706 19492 38708
tri 19492 38706 19494 38708 sw
tri 19250 38662 19294 38706 ne
rect 19294 38662 19494 38706
tri 19494 38662 19538 38706 sw
rect 70813 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19294 38620 19336 38662 ne
rect 19336 38620 19538 38662
tri 19336 38574 19382 38620 ne
rect 19382 38574 19458 38620
rect 19504 38604 19538 38620
tri 19538 38604 19596 38662 sw
rect 70813 38604 71000 38662
rect 19504 38574 19596 38604
tri 19382 38558 19398 38574 ne
rect 19398 38558 19596 38574
tri 19596 38558 19642 38604 sw
rect 70813 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
tri 19398 38500 19456 38558 ne
rect 19456 38500 19642 38558
tri 19642 38500 19700 38558 sw
rect 70813 38500 71000 38558
tri 19456 38488 19468 38500 ne
rect 19468 38488 19700 38500
tri 19700 38488 19712 38500 sw
tri 19468 38442 19514 38488 ne
rect 19514 38442 19590 38488
rect 19636 38454 19712 38488
tri 19712 38454 19746 38488 sw
rect 70813 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19746 38454
tri 19514 38396 19560 38442 ne
rect 19560 38396 19746 38442
tri 19746 38396 19804 38454 sw
rect 70813 38396 71000 38454
tri 19560 38356 19600 38396 ne
rect 19600 38356 19804 38396
tri 19804 38356 19844 38396 sw
tri 19600 38310 19646 38356 ne
rect 19646 38310 19722 38356
rect 19768 38350 19844 38356
tri 19844 38350 19850 38356 sw
rect 70813 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 19768 38310 19850 38350
tri 19850 38310 19890 38350 sw
tri 19646 38292 19664 38310 ne
rect 19664 38292 19890 38310
tri 19890 38292 19908 38310 sw
rect 70813 38292 71000 38350
tri 19664 38246 19710 38292 ne
rect 19710 38246 19908 38292
tri 19908 38246 19954 38292 sw
rect 70813 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
tri 19710 38224 19732 38246 ne
rect 19732 38240 19954 38246
tri 19954 38240 19960 38246 sw
rect 19732 38224 19960 38240
tri 19732 38178 19778 38224 ne
rect 19778 38178 19854 38224
rect 19900 38188 19960 38224
tri 19960 38188 20012 38240 sw
rect 70813 38188 71000 38246
rect 19900 38178 20012 38188
tri 19778 38142 19814 38178 ne
rect 19814 38142 20012 38178
tri 20012 38142 20058 38188 sw
rect 70813 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
tri 19814 38092 19864 38142 ne
rect 19864 38092 20058 38142
tri 20058 38092 20108 38142 sw
tri 19864 38046 19910 38092 ne
rect 19910 38046 19986 38092
rect 20032 38084 20108 38092
tri 20108 38084 20116 38092 sw
rect 70813 38084 71000 38142
rect 20032 38046 20116 38084
tri 20116 38046 20154 38084 sw
tri 19910 38038 19918 38046 ne
rect 19918 38038 20154 38046
tri 20154 38038 20162 38046 sw
rect 70813 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
tri 19918 37996 19960 38038 ne
rect 19960 37996 20162 38038
tri 19960 37980 19976 37996 ne
rect 19976 37980 20162 37996
tri 20162 37980 20220 38038 sw
rect 70813 37980 71000 38038
tri 19976 37960 19996 37980 ne
rect 19996 37960 20220 37980
tri 20220 37960 20240 37980 sw
tri 19996 37914 20042 37960 ne
rect 20042 37914 20118 37960
rect 20164 37934 20240 37960
tri 20240 37934 20266 37960 sw
rect 70813 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 20164 37914 20266 37934
tri 20266 37914 20286 37934 sw
tri 20042 37876 20080 37914 ne
rect 20080 37876 20286 37914
tri 20286 37876 20324 37914 sw
rect 70813 37876 71000 37934
tri 20080 37830 20126 37876 ne
rect 20126 37830 20324 37876
tri 20324 37830 20370 37876 sw
rect 70813 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
tri 20126 37828 20128 37830 ne
rect 20128 37828 20370 37830
tri 20370 37828 20372 37830 sw
tri 20128 37782 20174 37828 ne
rect 20174 37782 20250 37828
rect 20296 37782 20372 37828
tri 20174 37772 20184 37782 ne
rect 20184 37772 20372 37782
tri 20372 37772 20428 37828 sw
rect 70813 37772 71000 37830
tri 20184 37726 20230 37772 ne
rect 20230 37726 20428 37772
tri 20428 37726 20474 37772 sw
rect 70813 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
tri 20230 37696 20260 37726 ne
rect 20260 37696 20474 37726
tri 20474 37696 20504 37726 sw
tri 20260 37650 20306 37696 ne
rect 20306 37650 20382 37696
rect 20428 37668 20504 37696
tri 20504 37668 20532 37696 sw
rect 70813 37668 71000 37726
rect 20428 37650 20532 37668
tri 20532 37650 20550 37668 sw
tri 20306 37622 20334 37650 ne
rect 20334 37622 20550 37650
tri 20550 37622 20578 37650 sw
rect 70813 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20334 37564 20392 37622 ne
rect 20392 37564 20578 37622
tri 20578 37564 20636 37622 sw
rect 70813 37564 71000 37622
tri 20392 37518 20438 37564 ne
rect 20438 37518 20514 37564
rect 20560 37518 20636 37564
tri 20636 37518 20682 37564 sw
rect 70813 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
tri 20438 37460 20496 37518 ne
rect 20496 37460 20682 37518
tri 20682 37460 20740 37518 sw
rect 70813 37460 71000 37518
tri 20496 37432 20524 37460 ne
rect 20524 37432 20740 37460
tri 20740 37432 20768 37460 sw
tri 20524 37386 20570 37432 ne
rect 20570 37386 20646 37432
rect 20692 37414 20768 37432
tri 20768 37414 20786 37432 sw
rect 70813 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 20692 37386 20786 37414
tri 20570 37356 20600 37386 ne
rect 20600 37356 20786 37386
tri 20786 37356 20844 37414 sw
rect 70813 37356 71000 37414
tri 20600 37310 20646 37356 ne
rect 20646 37310 20844 37356
tri 20844 37310 20890 37356 sw
rect 70813 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
tri 20646 37300 20656 37310 ne
rect 20656 37300 20890 37310
tri 20890 37300 20900 37310 sw
tri 20656 37254 20702 37300 ne
rect 20702 37254 20778 37300
rect 20824 37254 20900 37300
tri 20900 37254 20946 37300 sw
tri 20702 37252 20704 37254 ne
rect 20704 37252 20946 37254
tri 20946 37252 20948 37254 sw
rect 70813 37252 71000 37310
tri 20704 37206 20750 37252 ne
rect 20750 37206 20948 37252
tri 20948 37206 20994 37252 sw
rect 70813 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
tri 20750 37168 20788 37206 ne
rect 20788 37168 20994 37206
tri 20788 37122 20834 37168 ne
rect 20834 37122 20910 37168
rect 20956 37148 20994 37168
tri 20994 37148 21052 37206 sw
rect 70813 37148 71000 37206
rect 20956 37122 21052 37148
tri 20834 37102 20854 37122 ne
rect 20854 37102 21052 37122
tri 21052 37102 21098 37148 sw
rect 70813 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20854 37044 20912 37102 ne
rect 20912 37044 21098 37102
tri 21098 37044 21156 37102 sw
rect 70813 37044 71000 37102
tri 20912 37036 20920 37044 ne
rect 20920 37036 21156 37044
tri 21156 37036 21164 37044 sw
tri 20920 36990 20966 37036 ne
rect 20966 36990 21042 37036
rect 21088 36998 21164 37036
tri 21164 36998 21202 37036 sw
rect 70813 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 21088 36990 21202 36998
tri 20966 36940 21016 36990 ne
rect 21016 36940 21202 36990
tri 21202 36940 21260 36998 sw
rect 70813 36940 71000 36998
tri 21016 36904 21052 36940 ne
rect 21052 36904 21260 36940
tri 21260 36904 21296 36940 sw
tri 21052 36858 21098 36904 ne
rect 21098 36858 21174 36904
rect 21220 36894 21296 36904
tri 21296 36894 21306 36904 sw
rect 70813 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 21220 36858 21306 36894
tri 21306 36858 21342 36894 sw
tri 21098 36836 21120 36858 ne
rect 21120 36836 21342 36858
tri 21342 36836 21364 36858 sw
rect 70813 36836 71000 36894
tri 21120 36790 21166 36836 ne
rect 21166 36790 21364 36836
tri 21364 36790 21410 36836 sw
rect 70813 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
tri 21166 36772 21184 36790 ne
rect 21184 36776 21410 36790
tri 21410 36776 21424 36790 sw
rect 21184 36772 21424 36776
tri 21184 36726 21230 36772 ne
rect 21230 36726 21306 36772
rect 21352 36732 21424 36772
tri 21424 36732 21468 36776 sw
rect 70813 36732 71000 36790
rect 21352 36726 21468 36732
tri 21230 36686 21270 36726 ne
rect 21270 36686 21468 36726
tri 21468 36686 21514 36732 sw
rect 70813 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
tri 21270 36640 21316 36686 ne
rect 21316 36640 21514 36686
tri 21514 36640 21560 36686 sw
tri 21316 36594 21362 36640 ne
rect 21362 36594 21438 36640
rect 21484 36628 21560 36640
tri 21560 36628 21572 36640 sw
rect 70813 36628 71000 36686
rect 21484 36594 21572 36628
tri 21572 36594 21606 36628 sw
tri 21362 36582 21374 36594 ne
rect 21374 36582 21606 36594
tri 21606 36582 21618 36594 sw
rect 70813 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21374 36532 21424 36582 ne
rect 21424 36532 21618 36582
tri 21424 36524 21432 36532 ne
rect 21432 36524 21618 36532
tri 21618 36524 21676 36582 sw
rect 70813 36524 71000 36582
tri 21432 36508 21448 36524 ne
rect 21448 36508 21676 36524
tri 21448 36462 21494 36508 ne
rect 21494 36462 21570 36508
rect 21616 36478 21676 36508
tri 21676 36478 21722 36524 sw
rect 70813 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 21616 36462 21722 36478
tri 21494 36420 21536 36462 ne
rect 21536 36420 21722 36462
tri 21722 36420 21780 36478 sw
rect 70813 36420 71000 36478
tri 21536 36376 21580 36420 ne
rect 21580 36376 21780 36420
tri 21780 36376 21824 36420 sw
tri 21580 36330 21626 36376 ne
rect 21626 36330 21702 36376
rect 21748 36374 21824 36376
tri 21824 36374 21826 36376 sw
rect 70813 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36330 21826 36374
tri 21626 36316 21640 36330 ne
rect 21640 36316 21826 36330
tri 21826 36316 21884 36374 sw
rect 70813 36316 71000 36374
tri 21640 36270 21686 36316 ne
rect 21686 36270 21884 36316
tri 21884 36270 21930 36316 sw
rect 70813 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
tri 21686 36244 21712 36270 ne
rect 21712 36244 21930 36270
tri 21930 36244 21956 36270 sw
tri 21712 36198 21758 36244 ne
rect 21758 36198 21834 36244
rect 21880 36212 21956 36244
tri 21956 36212 21988 36244 sw
rect 70813 36212 71000 36270
rect 21880 36198 21988 36212
tri 21988 36198 22002 36212 sw
tri 21758 36166 21790 36198 ne
rect 21790 36166 22002 36198
tri 22002 36166 22034 36198 sw
rect 70813 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21790 36112 21844 36166 ne
rect 21844 36112 22034 36166
tri 21844 36066 21890 36112 ne
rect 21890 36066 21966 36112
rect 22012 36108 22034 36112
tri 22034 36108 22092 36166 sw
rect 70813 36108 71000 36166
rect 22012 36066 22092 36108
tri 21890 36062 21894 36066 ne
rect 21894 36062 22092 36066
tri 22092 36062 22138 36108 sw
rect 70813 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
tri 21894 36004 21952 36062 ne
rect 21952 36004 22138 36062
tri 22138 36004 22196 36062 sw
rect 70813 36004 71000 36062
tri 21952 35980 21976 36004 ne
rect 21976 35980 22196 36004
tri 22196 35980 22220 36004 sw
tri 21976 35934 22022 35980 ne
rect 22022 35934 22098 35980
rect 22144 35958 22220 35980
tri 22220 35958 22242 35980 sw
rect 70813 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22144 35934 22242 35958
tri 22022 35900 22056 35934 ne
rect 22056 35900 22242 35934
tri 22242 35900 22300 35958 sw
rect 70813 35900 71000 35958
tri 22056 35854 22102 35900 ne
rect 22102 35854 22300 35900
tri 22300 35854 22346 35900 sw
rect 70813 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
tri 22102 35848 22108 35854 ne
rect 22108 35848 22346 35854
tri 22346 35848 22352 35854 sw
tri 22108 35802 22154 35848 ne
rect 22154 35802 22230 35848
rect 22276 35802 22352 35848
tri 22352 35802 22398 35848 sw
tri 22154 35796 22160 35802 ne
rect 22160 35796 22398 35802
tri 22398 35796 22404 35802 sw
rect 70813 35796 71000 35854
tri 22160 35750 22206 35796 ne
rect 22206 35750 22404 35796
tri 22404 35750 22450 35796 sw
rect 70813 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22206 35716 22240 35750 ne
rect 22240 35716 22450 35750
tri 22450 35716 22484 35750 sw
tri 22240 35670 22286 35716 ne
rect 22286 35670 22362 35716
rect 22408 35692 22484 35716
tri 22484 35692 22508 35716 sw
rect 70813 35692 71000 35750
rect 22408 35670 22508 35692
tri 22286 35646 22310 35670 ne
rect 22310 35646 22508 35670
tri 22508 35646 22554 35692 sw
rect 70813 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
tri 22310 35588 22368 35646 ne
rect 22368 35588 22554 35646
tri 22554 35588 22612 35646 sw
rect 70813 35588 71000 35646
tri 22368 35584 22372 35588 ne
rect 22372 35584 22612 35588
tri 22612 35584 22616 35588 sw
tri 22372 35538 22418 35584 ne
rect 22418 35538 22494 35584
rect 22540 35542 22616 35584
tri 22616 35542 22658 35584 sw
rect 70813 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 22540 35538 22658 35542
tri 22658 35538 22662 35542 sw
tri 22418 35484 22472 35538 ne
rect 22472 35484 22662 35538
tri 22662 35484 22716 35538 sw
rect 70813 35484 71000 35542
tri 22472 35452 22504 35484 ne
rect 22504 35452 22716 35484
tri 22504 35406 22550 35452 ne
rect 22550 35406 22626 35452
rect 22672 35438 22716 35452
tri 22716 35438 22762 35484 sw
rect 70813 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35406 22762 35438
tri 22550 35380 22576 35406 ne
rect 22576 35380 22762 35406
tri 22762 35380 22820 35438 sw
rect 70813 35380 71000 35438
tri 22576 35334 22622 35380 ne
rect 22622 35334 22820 35380
tri 22820 35334 22866 35380 sw
rect 70813 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
tri 22622 35320 22636 35334 ne
rect 22636 35320 22866 35334
tri 22866 35320 22880 35334 sw
tri 22636 35274 22682 35320 ne
rect 22682 35274 22758 35320
rect 22804 35276 22880 35320
tri 22880 35276 22924 35320 sw
rect 70813 35276 71000 35334
rect 22804 35274 22924 35276
tri 22682 35230 22726 35274 ne
rect 22726 35230 22924 35274
tri 22924 35230 22970 35276 sw
rect 70813 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22726 35188 22768 35230 ne
rect 22768 35188 22970 35230
tri 22970 35188 23012 35230 sw
tri 22768 35142 22814 35188 ne
rect 22814 35142 22890 35188
rect 22936 35172 23012 35188
tri 23012 35172 23028 35188 sw
rect 70813 35172 71000 35230
rect 22936 35142 23028 35172
tri 23028 35142 23058 35172 sw
tri 22814 35126 22830 35142 ne
rect 22830 35126 23058 35142
tri 23058 35126 23074 35142 sw
rect 70813 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
tri 22830 35068 22888 35126 ne
rect 22888 35068 23074 35126
tri 23074 35068 23132 35126 sw
rect 70813 35068 71000 35126
tri 22888 35056 22900 35068 ne
rect 22900 35056 23132 35068
tri 22900 35010 22946 35056 ne
rect 22946 35010 23022 35056
rect 23068 35022 23132 35056
tri 23132 35022 23178 35068 sw
rect 70813 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 23068 35010 23178 35022
tri 22946 34964 22992 35010 ne
rect 22992 34964 23178 35010
tri 23178 34964 23236 35022 sw
rect 70813 34964 71000 35022
tri 22992 34924 23032 34964 ne
rect 23032 34924 23236 34964
tri 23236 34924 23276 34964 sw
tri 23032 34878 23078 34924 ne
rect 23078 34878 23154 34924
rect 23200 34918 23276 34924
tri 23276 34918 23282 34924 sw
rect 70813 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34878 23282 34918
tri 23282 34878 23322 34918 sw
tri 23078 34860 23096 34878 ne
rect 23096 34860 23322 34878
tri 23322 34860 23340 34878 sw
rect 70813 34860 71000 34918
tri 23096 34824 23132 34860 ne
rect 23132 34824 23340 34860
tri 23132 34814 23142 34824 ne
rect 23142 34814 23340 34824
tri 23340 34814 23386 34860 sw
rect 70813 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
tri 23142 34792 23164 34814 ne
rect 23164 34792 23386 34814
tri 23164 34746 23210 34792 ne
rect 23210 34746 23286 34792
rect 23332 34756 23386 34792
tri 23386 34756 23444 34814 sw
rect 70813 34756 71000 34814
rect 23332 34746 23444 34756
tri 23210 34710 23246 34746 ne
rect 23246 34710 23444 34746
tri 23444 34710 23490 34756 sw
rect 70813 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23246 34660 23296 34710 ne
rect 23296 34660 23490 34710
tri 23490 34660 23540 34710 sw
tri 23296 34614 23342 34660 ne
rect 23342 34614 23418 34660
rect 23464 34652 23540 34660
tri 23540 34652 23548 34660 sw
rect 70813 34652 71000 34710
rect 23464 34614 23548 34652
tri 23342 34606 23350 34614 ne
rect 23350 34606 23548 34614
tri 23548 34606 23594 34652 sw
rect 70813 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
tri 23350 34548 23408 34606 ne
rect 23408 34548 23594 34606
tri 23594 34548 23652 34606 sw
rect 70813 34548 71000 34606
tri 23408 34528 23428 34548 ne
rect 23428 34528 23652 34548
tri 23652 34528 23672 34548 sw
tri 23428 34482 23474 34528 ne
rect 23474 34482 23550 34528
rect 23596 34502 23672 34528
tri 23672 34502 23698 34528 sw
rect 70813 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 23596 34482 23698 34502
tri 23698 34482 23718 34502 sw
tri 23474 34444 23512 34482 ne
rect 23512 34444 23718 34482
tri 23718 34444 23756 34482 sw
rect 70813 34444 71000 34502
tri 23512 34398 23558 34444 ne
rect 23558 34398 23756 34444
tri 23756 34398 23802 34444 sw
rect 70813 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
tri 23558 34396 23560 34398 ne
rect 23560 34396 23802 34398
tri 23560 34350 23606 34396 ne
rect 23606 34350 23682 34396
rect 23728 34350 23802 34396
tri 23606 34340 23616 34350 ne
rect 23616 34340 23802 34350
tri 23802 34340 23860 34398 sw
rect 70813 34340 71000 34398
tri 23616 34294 23662 34340 ne
rect 23662 34294 23860 34340
tri 23860 34294 23906 34340 sw
rect 70813 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23662 34264 23692 34294 ne
rect 23692 34264 23906 34294
tri 23906 34264 23936 34294 sw
tri 23692 34218 23738 34264 ne
rect 23738 34218 23814 34264
rect 23860 34236 23936 34264
tri 23936 34236 23964 34264 sw
rect 70813 34236 71000 34294
rect 23860 34218 23964 34236
tri 23738 34190 23766 34218 ne
rect 23766 34190 23964 34218
tri 23964 34190 24010 34236 sw
rect 70813 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
tri 23766 34132 23824 34190 ne
rect 23824 34132 24010 34190
tri 24010 34132 24068 34190 sw
rect 70813 34132 71000 34190
tri 23824 34086 23870 34132 ne
rect 23870 34086 23946 34132
rect 23992 34086 24068 34132
tri 24068 34086 24114 34132 sw
rect 70813 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
tri 23870 34028 23928 34086 ne
rect 23928 34028 24114 34086
tri 24114 34028 24172 34086 sw
rect 70813 34028 71000 34086
tri 23928 34000 23956 34028 ne
rect 23956 34000 24172 34028
tri 24172 34000 24200 34028 sw
tri 23956 33954 24002 34000 ne
rect 24002 33954 24078 34000
rect 24124 33982 24200 34000
tri 24200 33982 24218 34000 sw
rect 70813 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33954 24218 33982
tri 24002 33924 24032 33954 ne
rect 24032 33924 24218 33954
tri 24218 33924 24276 33982 sw
rect 70813 33924 71000 33982
tri 24032 33878 24078 33924 ne
rect 24078 33878 24276 33924
tri 24276 33878 24322 33924 sw
rect 70813 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
tri 24078 33868 24088 33878 ne
rect 24088 33868 24322 33878
tri 24322 33868 24332 33878 sw
tri 24088 33822 24134 33868 ne
rect 24134 33822 24210 33868
rect 24256 33822 24332 33868
tri 24332 33822 24378 33868 sw
tri 24134 33820 24136 33822 ne
rect 24136 33820 24378 33822
tri 24378 33820 24380 33822 sw
rect 70813 33820 71000 33878
tri 24136 33774 24182 33820 ne
rect 24182 33774 24380 33820
tri 24380 33774 24426 33820 sw
rect 70813 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24182 33736 24220 33774 ne
rect 24220 33736 24426 33774
tri 24220 33690 24266 33736 ne
rect 24266 33690 24342 33736
rect 24388 33716 24426 33736
tri 24426 33716 24484 33774 sw
rect 70813 33716 71000 33774
rect 24388 33690 24484 33716
tri 24266 33670 24286 33690 ne
rect 24286 33670 24484 33690
tri 24484 33670 24530 33716 sw
rect 70813 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
tri 24286 33612 24344 33670 ne
rect 24344 33612 24530 33670
tri 24530 33612 24588 33670 sw
rect 70813 33612 71000 33670
tri 24344 33604 24352 33612 ne
rect 24352 33604 24588 33612
tri 24588 33604 24596 33612 sw
tri 24352 33558 24398 33604 ne
rect 24398 33558 24474 33604
rect 24520 33566 24596 33604
tri 24596 33566 24634 33604 sw
rect 70813 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 24520 33558 24634 33566
tri 24398 33508 24448 33558 ne
rect 24448 33508 24634 33558
tri 24634 33508 24692 33566 sw
rect 70813 33508 71000 33566
tri 24448 33472 24484 33508 ne
rect 24484 33472 24692 33508
tri 24692 33472 24728 33508 sw
tri 24484 33426 24530 33472 ne
rect 24530 33426 24606 33472
rect 24652 33462 24728 33472
tri 24728 33462 24738 33472 sw
rect 70813 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24652 33426 24738 33462
tri 24738 33426 24774 33462 sw
tri 24530 33404 24552 33426 ne
rect 24552 33404 24774 33426
tri 24774 33404 24796 33426 sw
rect 70813 33404 71000 33462
tri 24552 33358 24598 33404 ne
rect 24598 33358 24796 33404
tri 24796 33358 24842 33404 sw
rect 70813 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
tri 24598 33340 24616 33358 ne
rect 24616 33340 24842 33358
tri 24616 33294 24662 33340 ne
rect 24662 33294 24738 33340
rect 24784 33300 24842 33340
tri 24842 33300 24900 33358 sw
rect 70813 33300 71000 33358
rect 24784 33294 24900 33300
tri 24662 33254 24702 33294 ne
rect 24702 33254 24900 33294
tri 24900 33254 24946 33300 sw
rect 70813 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24702 33208 24748 33254 ne
rect 24748 33208 24946 33254
tri 24946 33208 24992 33254 sw
tri 24748 33162 24794 33208 ne
rect 24794 33162 24870 33208
rect 24916 33196 24992 33208
tri 24992 33196 25004 33208 sw
rect 70813 33196 71000 33254
rect 24916 33162 25004 33196
tri 25004 33162 25038 33196 sw
tri 24794 33150 24806 33162 ne
rect 24806 33150 25038 33162
tri 25038 33150 25050 33162 sw
rect 70813 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
tri 24806 33116 24840 33150 ne
rect 24840 33116 25050 33150
tri 24840 33092 24864 33116 ne
rect 24864 33092 25050 33116
tri 25050 33092 25108 33150 sw
rect 70813 33092 71000 33150
tri 24864 33076 24880 33092 ne
rect 24880 33076 25108 33092
tri 24880 33030 24926 33076 ne
rect 24926 33030 25002 33076
rect 25048 33046 25108 33076
tri 25108 33046 25154 33092 sw
rect 70813 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 25048 33030 25154 33046
tri 24926 32988 24968 33030 ne
rect 24968 32988 25154 33030
tri 25154 32988 25212 33046 sw
rect 70813 32988 71000 33046
tri 24968 32944 25012 32988 ne
rect 25012 32944 25212 32988
tri 25212 32944 25256 32988 sw
tri 25012 32898 25058 32944 ne
rect 25058 32898 25134 32944
rect 25180 32942 25256 32944
tri 25256 32942 25258 32944 sw
rect 70813 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32898 25258 32942
tri 25058 32884 25072 32898 ne
rect 25072 32884 25258 32898
tri 25258 32884 25316 32942 sw
rect 70813 32884 71000 32942
tri 25072 32838 25118 32884 ne
rect 25118 32838 25316 32884
tri 25316 32838 25362 32884 sw
rect 70813 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
tri 25118 32812 25144 32838 ne
rect 25144 32812 25362 32838
tri 25362 32812 25388 32838 sw
tri 25144 32766 25190 32812 ne
rect 25190 32766 25266 32812
rect 25312 32780 25388 32812
tri 25388 32780 25420 32812 sw
rect 70813 32780 71000 32838
rect 25312 32766 25420 32780
tri 25420 32766 25434 32780 sw
tri 25190 32734 25222 32766 ne
rect 25222 32734 25434 32766
tri 25434 32734 25466 32766 sw
rect 70813 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25222 32680 25276 32734 ne
rect 25276 32680 25466 32734
tri 25276 32634 25322 32680 ne
rect 25322 32634 25398 32680
rect 25444 32676 25466 32680
tri 25466 32676 25524 32734 sw
rect 70813 32676 71000 32734
rect 25444 32634 25524 32676
tri 25322 32630 25326 32634 ne
rect 25326 32630 25524 32634
tri 25524 32630 25570 32676 sw
rect 70813 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25326 32572 25384 32630 ne
rect 25384 32572 25570 32630
tri 25570 32572 25628 32630 sw
rect 70813 32572 71000 32630
tri 25384 32548 25408 32572 ne
rect 25408 32548 25628 32572
tri 25628 32548 25652 32572 sw
tri 25408 32502 25454 32548 ne
rect 25454 32502 25530 32548
rect 25576 32526 25652 32548
tri 25652 32526 25674 32548 sw
rect 70813 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 25576 32502 25674 32526
tri 25454 32468 25488 32502 ne
rect 25488 32468 25674 32502
tri 25674 32468 25732 32526 sw
rect 70813 32468 71000 32526
tri 25488 32422 25534 32468 ne
rect 25534 32422 25732 32468
tri 25732 32422 25778 32468 sw
rect 70813 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
tri 25534 32416 25540 32422 ne
rect 25540 32416 25778 32422
tri 25778 32416 25784 32422 sw
tri 25540 32370 25586 32416 ne
rect 25586 32370 25662 32416
rect 25708 32370 25784 32416
tri 25784 32370 25830 32416 sw
tri 25586 32364 25592 32370 ne
rect 25592 32364 25830 32370
tri 25830 32364 25836 32370 sw
rect 70813 32364 71000 32422
tri 25592 32318 25638 32364 ne
rect 25638 32318 25836 32364
tri 25836 32318 25882 32364 sw
rect 70813 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
tri 25638 32284 25672 32318 ne
rect 25672 32284 25882 32318
tri 25882 32284 25916 32318 sw
tri 25672 32238 25718 32284 ne
rect 25718 32238 25794 32284
rect 25840 32260 25916 32284
tri 25916 32260 25940 32284 sw
rect 70813 32260 71000 32318
rect 25840 32238 25940 32260
tri 25718 32214 25742 32238 ne
rect 25742 32214 25940 32238
tri 25940 32214 25986 32260 sw
rect 70813 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25742 32156 25800 32214 ne
rect 25800 32156 25986 32214
tri 25986 32156 26044 32214 sw
rect 70813 32156 71000 32214
tri 25800 32152 25804 32156 ne
rect 25804 32152 26044 32156
tri 26044 32152 26048 32156 sw
tri 25804 32106 25850 32152 ne
rect 25850 32106 25926 32152
rect 25972 32110 26048 32152
tri 26048 32110 26090 32152 sw
rect 70813 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 25972 32106 26090 32110
tri 26090 32106 26094 32110 sw
tri 25850 32052 25904 32106 ne
rect 25904 32052 26094 32106
tri 26094 32052 26148 32106 sw
rect 70813 32052 71000 32110
tri 25904 32020 25936 32052 ne
rect 25936 32020 26148 32052
tri 25936 31974 25982 32020 ne
rect 25982 31974 26058 32020
rect 26104 32006 26148 32020
tri 26148 32006 26194 32052 sw
rect 70813 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 26104 31974 26194 32006
tri 25982 31948 26008 31974 ne
rect 26008 31948 26194 31974
tri 26194 31948 26252 32006 sw
rect 70813 31948 71000 32006
tri 26008 31902 26054 31948 ne
rect 26054 31902 26252 31948
tri 26252 31902 26298 31948 sw
rect 70813 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
tri 26054 31888 26068 31902 ne
rect 26068 31888 26298 31902
tri 26298 31888 26312 31902 sw
tri 26068 31842 26114 31888 ne
rect 26114 31842 26190 31888
rect 26236 31844 26312 31888
tri 26312 31844 26356 31888 sw
rect 70813 31844 71000 31902
rect 26236 31842 26356 31844
tri 26114 31798 26158 31842 ne
rect 26158 31798 26356 31842
tri 26356 31798 26402 31844 sw
rect 70813 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
tri 26158 31756 26200 31798 ne
rect 26200 31756 26402 31798
tri 26402 31756 26444 31798 sw
tri 26200 31710 26246 31756 ne
rect 26246 31710 26322 31756
rect 26368 31740 26444 31756
tri 26444 31740 26460 31756 sw
rect 70813 31740 71000 31798
rect 26368 31710 26460 31740
tri 26460 31710 26490 31740 sw
tri 26246 31694 26262 31710 ne
rect 26262 31694 26490 31710
tri 26490 31694 26506 31710 sw
rect 70813 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
tri 26262 31636 26320 31694 ne
rect 26320 31636 26506 31694
tri 26506 31636 26564 31694 sw
rect 70813 31636 71000 31694
tri 26320 31624 26332 31636 ne
rect 26332 31624 26564 31636
tri 26332 31578 26378 31624 ne
rect 26378 31578 26454 31624
rect 26500 31590 26564 31624
tri 26564 31590 26610 31636 sw
rect 70813 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 26500 31578 26610 31590
tri 26378 31532 26424 31578 ne
rect 26424 31532 26610 31578
tri 26610 31532 26668 31590 sw
rect 70813 31532 71000 31590
tri 26424 31492 26464 31532 ne
rect 26464 31492 26668 31532
tri 26668 31492 26708 31532 sw
tri 26464 31446 26510 31492 ne
rect 26510 31446 26586 31492
rect 26632 31486 26708 31492
tri 26708 31486 26714 31492 sw
rect 70813 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31446 26714 31486
tri 26714 31446 26754 31486 sw
tri 26510 31428 26528 31446 ne
rect 26528 31428 26754 31446
tri 26754 31428 26772 31446 sw
rect 70813 31428 71000 31486
tri 26528 31408 26548 31428 ne
rect 26548 31408 26772 31428
tri 26548 31382 26574 31408 ne
rect 26574 31382 26772 31408
tri 26772 31382 26818 31428 sw
rect 70813 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
tri 26574 31360 26596 31382 ne
rect 26596 31360 26818 31382
tri 26596 31314 26642 31360 ne
rect 26642 31314 26718 31360
rect 26764 31324 26818 31360
tri 26818 31324 26876 31382 sw
rect 70813 31324 71000 31382
rect 26764 31314 26876 31324
tri 26642 31278 26678 31314 ne
rect 26678 31278 26876 31314
tri 26876 31278 26922 31324 sw
rect 70813 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
tri 26678 31228 26728 31278 ne
rect 26728 31228 26922 31278
tri 26922 31228 26972 31278 sw
tri 26728 31182 26774 31228 ne
rect 26774 31182 26850 31228
rect 26896 31220 26972 31228
tri 26972 31220 26980 31228 sw
rect 70813 31220 71000 31278
rect 26896 31182 26980 31220
tri 26774 31174 26782 31182 ne
rect 26782 31174 26980 31182
tri 26980 31174 27026 31220 sw
rect 70813 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
tri 26782 31116 26840 31174 ne
rect 26840 31116 27026 31174
tri 27026 31116 27084 31174 sw
rect 70813 31116 71000 31174
tri 26840 31096 26860 31116 ne
rect 26860 31096 27084 31116
tri 27084 31096 27104 31116 sw
tri 26860 31050 26906 31096 ne
rect 26906 31050 26982 31096
rect 27028 31070 27104 31096
tri 27104 31070 27130 31096 sw
rect 70813 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 27028 31050 27130 31070
tri 27130 31050 27150 31070 sw
tri 26906 31012 26944 31050 ne
rect 26944 31012 27150 31050
tri 27150 31012 27188 31050 sw
rect 70813 31012 71000 31070
tri 26944 30966 26990 31012 ne
rect 26990 30966 27188 31012
tri 27188 30966 27234 31012 sw
rect 70813 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
tri 26990 30964 26992 30966 ne
rect 26992 30964 27234 30966
tri 26992 30918 27038 30964 ne
rect 27038 30918 27114 30964
rect 27160 30918 27234 30964
tri 27038 30908 27048 30918 ne
rect 27048 30908 27234 30918
tri 27234 30908 27292 30966 sw
rect 70813 30908 71000 30966
tri 27048 30862 27094 30908 ne
rect 27094 30862 27292 30908
tri 27292 30862 27338 30908 sw
rect 70813 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
tri 27094 30832 27124 30862 ne
rect 27124 30832 27338 30862
tri 27338 30832 27368 30862 sw
tri 27124 30786 27170 30832 ne
rect 27170 30786 27246 30832
rect 27292 30804 27368 30832
tri 27368 30804 27396 30832 sw
rect 70813 30804 71000 30862
rect 27292 30786 27396 30804
tri 27170 30758 27198 30786 ne
rect 27198 30758 27396 30786
tri 27396 30758 27442 30804 sw
rect 70813 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27198 30700 27256 30758 ne
rect 27256 30700 27442 30758
tri 27442 30700 27500 30758 sw
rect 70813 30700 71000 30758
tri 27256 30654 27302 30700 ne
rect 27302 30654 27378 30700
rect 27424 30654 27500 30700
tri 27500 30654 27546 30700 sw
rect 70813 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
tri 27302 30596 27360 30654 ne
rect 27360 30596 27546 30654
tri 27546 30596 27604 30654 sw
rect 70813 30596 71000 30654
tri 27360 30568 27388 30596 ne
rect 27388 30568 27604 30596
tri 27604 30568 27632 30596 sw
tri 27388 30522 27434 30568 ne
rect 27434 30522 27510 30568
rect 27556 30550 27632 30568
tri 27632 30550 27650 30568 sw
rect 70813 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30522 27650 30550
tri 27434 30492 27464 30522 ne
rect 27464 30492 27650 30522
tri 27650 30492 27708 30550 sw
rect 70813 30492 71000 30550
tri 27464 30446 27510 30492 ne
rect 27510 30446 27708 30492
tri 27708 30446 27754 30492 sw
rect 70813 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
tri 27510 30436 27520 30446 ne
rect 27520 30436 27754 30446
tri 27754 30436 27764 30446 sw
tri 27520 30390 27566 30436 ne
rect 27566 30390 27642 30436
rect 27688 30390 27764 30436
tri 27764 30390 27810 30436 sw
tri 27566 30388 27568 30390 ne
rect 27568 30388 27810 30390
tri 27810 30388 27812 30390 sw
rect 70813 30388 71000 30446
tri 27568 30342 27614 30388 ne
rect 27614 30342 27812 30388
tri 27812 30342 27858 30388 sw
rect 70813 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27614 30304 27652 30342 ne
rect 27652 30304 27858 30342
tri 27652 30258 27698 30304 ne
rect 27698 30258 27774 30304
rect 27820 30284 27858 30304
tri 27858 30284 27916 30342 sw
rect 70813 30284 71000 30342
rect 27820 30258 27916 30284
tri 27698 30238 27718 30258 ne
rect 27718 30238 27916 30258
tri 27916 30238 27962 30284 sw
rect 70813 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27718 30180 27776 30238 ne
rect 27776 30180 27962 30238
tri 27962 30180 28020 30238 sw
rect 70813 30180 71000 30238
tri 27776 30172 27784 30180 ne
rect 27784 30172 28020 30180
tri 28020 30172 28028 30180 sw
tri 27784 30126 27830 30172 ne
rect 27830 30126 27906 30172
rect 27952 30134 28028 30172
tri 28028 30134 28066 30172 sw
rect 70813 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 27952 30126 28066 30134
tri 27830 30076 27880 30126 ne
rect 27880 30076 28066 30126
tri 28066 30076 28124 30134 sw
rect 70813 30076 71000 30134
tri 27880 30040 27916 30076 ne
rect 27916 30040 28124 30076
tri 28124 30040 28160 30076 sw
tri 27916 29994 27962 30040 ne
rect 27962 29994 28038 30040
rect 28084 30030 28160 30040
tri 28160 30030 28170 30040 sw
rect 70813 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 29994 28170 30030
tri 28170 29994 28206 30030 sw
tri 27962 29972 27984 29994 ne
rect 27984 29972 28206 29994
tri 28206 29972 28228 29994 sw
rect 70813 29972 71000 30030
tri 27984 29926 28030 29972 ne
rect 28030 29926 28228 29972
tri 28228 29926 28274 29972 sw
rect 70813 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
tri 28030 29908 28048 29926 ne
rect 28048 29908 28274 29926
tri 28048 29862 28094 29908 ne
rect 28094 29862 28170 29908
rect 28216 29868 28274 29908
tri 28274 29868 28332 29926 sw
rect 70813 29868 71000 29926
rect 28216 29862 28332 29868
tri 28094 29822 28134 29862 ne
rect 28134 29822 28332 29862
tri 28332 29822 28378 29868 sw
rect 70813 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
tri 28134 29776 28180 29822 ne
rect 28180 29776 28378 29822
tri 28378 29776 28424 29822 sw
tri 28180 29730 28226 29776 ne
rect 28226 29730 28302 29776
rect 28348 29764 28424 29776
tri 28424 29764 28436 29776 sw
rect 70813 29764 71000 29822
rect 28348 29730 28436 29764
tri 28436 29730 28470 29764 sw
tri 28226 29718 28238 29730 ne
rect 28238 29718 28470 29730
tri 28470 29718 28482 29730 sw
rect 70813 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
tri 28238 29700 28256 29718 ne
rect 28256 29700 28482 29718
tri 28256 29660 28296 29700 ne
rect 28296 29660 28482 29700
tri 28482 29660 28540 29718 sw
rect 70813 29660 71000 29718
tri 28296 29644 28312 29660 ne
rect 28312 29644 28540 29660
tri 28312 29598 28358 29644 ne
rect 28358 29598 28434 29644
rect 28480 29614 28540 29644
tri 28540 29614 28586 29660 sw
rect 70813 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 28480 29598 28586 29614
tri 28358 29556 28400 29598 ne
rect 28400 29556 28586 29598
tri 28586 29556 28644 29614 sw
rect 70813 29556 71000 29614
tri 28400 29512 28444 29556 ne
rect 28444 29512 28644 29556
tri 28644 29512 28688 29556 sw
tri 28444 29466 28490 29512 ne
rect 28490 29466 28566 29512
rect 28612 29510 28688 29512
tri 28688 29510 28690 29512 sw
rect 70813 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29466 28690 29510
tri 28490 29452 28504 29466 ne
rect 28504 29452 28690 29466
tri 28690 29452 28748 29510 sw
rect 70813 29452 71000 29510
tri 28504 29406 28550 29452 ne
rect 28550 29406 28748 29452
tri 28748 29406 28794 29452 sw
rect 70813 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28550 29380 28576 29406 ne
rect 28576 29380 28794 29406
tri 28794 29380 28820 29406 sw
tri 28576 29334 28622 29380 ne
rect 28622 29334 28698 29380
rect 28744 29348 28820 29380
tri 28820 29348 28852 29380 sw
rect 70813 29348 71000 29406
rect 28744 29334 28852 29348
tri 28852 29334 28866 29348 sw
tri 28622 29302 28654 29334 ne
rect 28654 29302 28866 29334
tri 28866 29302 28898 29334 sw
rect 70813 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28654 29248 28708 29302 ne
rect 28708 29248 28898 29302
tri 28708 29202 28754 29248 ne
rect 28754 29202 28830 29248
rect 28876 29244 28898 29248
tri 28898 29244 28956 29302 sw
rect 70813 29244 71000 29302
rect 28876 29202 28956 29244
tri 28754 29198 28758 29202 ne
rect 28758 29198 28956 29202
tri 28956 29198 29002 29244 sw
rect 70813 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
tri 28758 29140 28816 29198 ne
rect 28816 29140 29002 29198
tri 29002 29140 29060 29198 sw
rect 70813 29140 71000 29198
tri 28816 29116 28840 29140 ne
rect 28840 29116 29060 29140
tri 29060 29116 29084 29140 sw
tri 28840 29070 28886 29116 ne
rect 28886 29070 28962 29116
rect 29008 29094 29084 29116
tri 29084 29094 29106 29116 sw
rect 70813 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 29008 29070 29106 29094
tri 28886 29036 28920 29070 ne
rect 28920 29036 29106 29070
tri 29106 29036 29164 29094 sw
rect 70813 29036 71000 29094
tri 28920 28990 28966 29036 ne
rect 28966 28990 29164 29036
tri 29164 28990 29210 29036 sw
rect 70813 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
tri 28966 28984 28972 28990 ne
rect 28972 28984 29210 28990
tri 29210 28984 29216 28990 sw
tri 28972 28938 29018 28984 ne
rect 29018 28938 29094 28984
rect 29140 28938 29216 28984
tri 29216 28938 29262 28984 sw
tri 29018 28932 29024 28938 ne
rect 29024 28932 29262 28938
tri 29262 28932 29268 28938 sw
rect 70813 28932 71000 28990
tri 29024 28886 29070 28932 ne
rect 29070 28886 29268 28932
tri 29268 28886 29314 28932 sw
rect 70813 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29070 28852 29104 28886 ne
rect 29104 28852 29314 28886
tri 29314 28852 29348 28886 sw
tri 29104 28806 29150 28852 ne
rect 29150 28806 29226 28852
rect 29272 28828 29348 28852
tri 29348 28828 29372 28852 sw
rect 70813 28828 71000 28886
rect 29272 28806 29372 28828
tri 29150 28782 29174 28806 ne
rect 29174 28782 29372 28806
tri 29372 28782 29418 28828 sw
rect 70813 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
tri 29174 28724 29232 28782 ne
rect 29232 28724 29418 28782
tri 29418 28724 29476 28782 sw
rect 70813 28724 71000 28782
tri 29232 28720 29236 28724 ne
rect 29236 28720 29476 28724
tri 29476 28720 29480 28724 sw
tri 29236 28674 29282 28720 ne
rect 29282 28674 29358 28720
rect 29404 28678 29480 28720
tri 29480 28678 29522 28720 sw
rect 70813 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 29404 28674 29522 28678
tri 29522 28674 29526 28678 sw
tri 29282 28620 29336 28674 ne
rect 29336 28620 29526 28674
tri 29526 28620 29580 28674 sw
rect 70813 28620 71000 28678
tri 29336 28588 29368 28620 ne
rect 29368 28588 29580 28620
tri 29368 28542 29414 28588 ne
rect 29414 28542 29490 28588
rect 29536 28574 29580 28588
tri 29580 28574 29626 28620 sw
rect 70813 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28542 29626 28574
tri 29414 28516 29440 28542 ne
rect 29440 28516 29626 28542
tri 29626 28516 29684 28574 sw
rect 70813 28516 71000 28574
tri 29440 28470 29486 28516 ne
rect 29486 28470 29684 28516
tri 29684 28470 29730 28516 sw
rect 70813 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
tri 29486 28456 29500 28470 ne
rect 29500 28456 29730 28470
tri 29730 28456 29744 28470 sw
tri 29500 28410 29546 28456 ne
rect 29546 28410 29622 28456
rect 29668 28412 29744 28456
tri 29744 28412 29788 28456 sw
rect 70813 28412 71000 28470
rect 29668 28410 29788 28412
tri 29546 28366 29590 28410 ne
rect 29590 28366 29788 28410
tri 29788 28366 29834 28412 sw
rect 70813 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29590 28324 29632 28366 ne
rect 29632 28324 29834 28366
tri 29834 28324 29876 28366 sw
tri 29632 28278 29678 28324 ne
rect 29678 28278 29754 28324
rect 29800 28308 29876 28324
tri 29876 28308 29892 28324 sw
rect 70813 28308 71000 28366
rect 29800 28278 29892 28308
tri 29892 28278 29922 28308 sw
tri 29678 28262 29694 28278 ne
rect 29694 28262 29922 28278
tri 29922 28262 29938 28278 sw
rect 70813 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
tri 29694 28204 29752 28262 ne
rect 29752 28204 29938 28262
tri 29938 28204 29996 28262 sw
rect 70813 28204 71000 28262
tri 29752 28192 29764 28204 ne
rect 29764 28192 29996 28204
tri 29764 28146 29810 28192 ne
rect 29810 28146 29886 28192
rect 29932 28158 29996 28192
tri 29996 28158 30042 28204 sw
rect 70813 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 29932 28146 30042 28158
tri 29810 28100 29856 28146 ne
rect 29856 28100 30042 28146
tri 30042 28100 30100 28158 sw
rect 70813 28100 71000 28158
tri 29856 28060 29896 28100 ne
rect 29896 28060 30100 28100
tri 30100 28060 30140 28100 sw
tri 29896 28014 29942 28060 ne
rect 29942 28014 30018 28060
rect 30064 28054 30140 28060
tri 30140 28054 30146 28060 sw
rect 70813 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28014 30146 28054
tri 30146 28014 30186 28054 sw
tri 29942 27996 29960 28014 ne
rect 29960 27996 30186 28014
tri 30186 27996 30204 28014 sw
rect 70813 27996 71000 28054
tri 29960 27992 29964 27996 ne
rect 29964 27992 30204 27996
tri 29964 27950 30006 27992 ne
rect 30006 27950 30204 27992
tri 30204 27950 30250 27996 sw
rect 70813 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
tri 30006 27928 30028 27950 ne
rect 30028 27928 30250 27950
tri 30028 27882 30074 27928 ne
rect 30074 27882 30150 27928
rect 30196 27892 30250 27928
tri 30250 27892 30308 27950 sw
rect 70813 27892 71000 27950
rect 30196 27882 30308 27892
tri 30074 27846 30110 27882 ne
rect 30110 27846 30308 27882
tri 30308 27846 30354 27892 sw
rect 70813 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30110 27796 30160 27846 ne
rect 30160 27796 30354 27846
tri 30354 27796 30404 27846 sw
tri 30160 27750 30206 27796 ne
rect 30206 27750 30282 27796
rect 30328 27788 30404 27796
tri 30404 27788 30412 27796 sw
rect 70813 27788 71000 27846
rect 30328 27750 30412 27788
tri 30206 27742 30214 27750 ne
rect 30214 27742 30412 27750
tri 30412 27742 30458 27788 sw
rect 70813 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
tri 30214 27684 30272 27742 ne
rect 30272 27684 30458 27742
tri 30458 27684 30516 27742 sw
rect 70813 27684 71000 27742
tri 30272 27664 30292 27684 ne
rect 30292 27664 30516 27684
tri 30516 27664 30536 27684 sw
tri 30292 27618 30338 27664 ne
rect 30338 27618 30414 27664
rect 30460 27638 30536 27664
tri 30536 27638 30562 27664 sw
rect 70813 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30460 27618 30562 27638
tri 30562 27618 30582 27638 sw
tri 30338 27580 30376 27618 ne
rect 30376 27580 30582 27618
tri 30582 27580 30620 27618 sw
rect 70813 27580 71000 27638
tri 30376 27534 30422 27580 ne
rect 30422 27534 30620 27580
tri 30620 27534 30666 27580 sw
rect 70813 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
tri 30422 27532 30424 27534 ne
rect 30424 27532 30666 27534
tri 30424 27486 30470 27532 ne
rect 30470 27486 30546 27532
rect 30592 27486 30666 27532
tri 30470 27476 30480 27486 ne
rect 30480 27476 30666 27486
tri 30666 27476 30724 27534 sw
rect 70813 27476 71000 27534
tri 30480 27430 30526 27476 ne
rect 30526 27430 30724 27476
tri 30724 27430 30770 27476 sw
rect 70813 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30526 27400 30556 27430 ne
rect 30556 27400 30770 27430
tri 30770 27400 30800 27430 sw
tri 30556 27354 30602 27400 ne
rect 30602 27354 30678 27400
rect 30724 27372 30800 27400
tri 30800 27372 30828 27400 sw
rect 70813 27372 71000 27430
rect 30724 27354 30828 27372
tri 30602 27326 30630 27354 ne
rect 30630 27326 30828 27354
tri 30828 27326 30874 27372 sw
rect 70813 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
tri 30630 27268 30688 27326 ne
rect 30688 27268 30874 27326
tri 30874 27268 30932 27326 sw
rect 70813 27268 71000 27326
tri 30688 27222 30734 27268 ne
rect 30734 27222 30810 27268
rect 30856 27222 30932 27268
tri 30932 27222 30978 27268 sw
rect 70813 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30734 27164 30792 27222 ne
rect 30792 27164 30978 27222
tri 30978 27164 31036 27222 sw
rect 70813 27164 71000 27222
tri 30792 27136 30820 27164 ne
rect 30820 27136 31036 27164
tri 31036 27136 31064 27164 sw
tri 30820 27090 30866 27136 ne
rect 30866 27090 30942 27136
rect 30988 27118 31064 27136
tri 31064 27118 31082 27136 sw
rect 70813 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 30988 27090 31082 27118
tri 30866 27060 30896 27090 ne
rect 30896 27060 31082 27090
tri 31082 27060 31140 27118 sw
rect 70813 27060 71000 27118
tri 30896 27014 30942 27060 ne
rect 30942 27014 31140 27060
tri 31140 27014 31186 27060 sw
rect 70813 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
tri 30942 27004 30952 27014 ne
rect 30952 27004 31186 27014
tri 31186 27004 31196 27014 sw
tri 30952 26958 30998 27004 ne
rect 30998 26958 31074 27004
rect 31120 26958 31196 27004
tri 31196 26958 31242 27004 sw
tri 30998 26956 31000 26958 ne
rect 31000 26956 31242 26958
tri 31242 26956 31244 26958 sw
rect 70813 26956 71000 27014
tri 31000 26910 31046 26956 ne
rect 31046 26910 31244 26956
tri 31244 26910 31290 26956 sw
rect 70813 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31046 26872 31084 26910 ne
rect 31084 26872 31290 26910
tri 31084 26826 31130 26872 ne
rect 31130 26826 31206 26872
rect 31252 26852 31290 26872
tri 31290 26852 31348 26910 sw
rect 70813 26852 71000 26910
rect 31252 26826 31348 26852
tri 31130 26806 31150 26826 ne
rect 31150 26806 31348 26826
tri 31348 26806 31394 26852 sw
rect 70813 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
tri 31150 26748 31208 26806 ne
rect 31208 26748 31394 26806
tri 31394 26748 31452 26806 sw
rect 70813 26748 71000 26806
tri 31208 26740 31216 26748 ne
rect 31216 26740 31452 26748
tri 31452 26740 31460 26748 sw
tri 31216 26694 31262 26740 ne
rect 31262 26694 31338 26740
rect 31384 26702 31460 26740
tri 31460 26702 31498 26740 sw
rect 70813 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 31384 26694 31498 26702
tri 31262 26644 31312 26694 ne
rect 31312 26644 31498 26694
tri 31498 26644 31556 26702 sw
rect 70813 26644 71000 26702
tri 31312 26608 31348 26644 ne
rect 31348 26608 31556 26644
tri 31556 26608 31592 26644 sw
tri 31348 26562 31394 26608 ne
rect 31394 26562 31470 26608
rect 31516 26598 31592 26608
tri 31592 26598 31602 26608 sw
rect 70813 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 31516 26562 31602 26598
tri 31602 26562 31638 26598 sw
tri 31394 26540 31416 26562 ne
rect 31416 26540 31638 26562
tri 31638 26540 31660 26562 sw
rect 70813 26540 71000 26598
tri 31416 26494 31462 26540 ne
rect 31462 26494 31660 26540
tri 31660 26494 31706 26540 sw
rect 70813 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
tri 31462 26476 31480 26494 ne
rect 31480 26476 31706 26494
tri 31480 26430 31526 26476 ne
rect 31526 26430 31602 26476
rect 31648 26436 31706 26476
tri 31706 26436 31764 26494 sw
rect 70813 26436 71000 26494
rect 31648 26430 31764 26436
tri 31526 26390 31566 26430 ne
rect 31566 26390 31764 26430
tri 31764 26390 31810 26436 sw
rect 70813 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31566 26344 31612 26390 ne
rect 31612 26344 31810 26390
tri 31810 26344 31856 26390 sw
tri 31612 26298 31658 26344 ne
rect 31658 26298 31734 26344
rect 31780 26332 31856 26344
tri 31856 26332 31868 26344 sw
rect 70813 26332 71000 26390
rect 31780 26298 31868 26332
tri 31868 26298 31902 26332 sw
tri 31658 26286 31670 26298 ne
rect 31670 26286 31902 26298
tri 31902 26286 31914 26298 sw
rect 70813 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31670 26284 31672 26286 ne
rect 31672 26284 31914 26286
tri 31672 26228 31728 26284 ne
rect 31728 26228 31914 26284
tri 31914 26228 31972 26286 sw
rect 70813 26228 71000 26286
tri 31728 26212 31744 26228 ne
rect 31744 26212 31972 26228
tri 31744 26166 31790 26212 ne
rect 31790 26166 31866 26212
rect 31912 26182 31972 26212
tri 31972 26182 32018 26228 sw
rect 70813 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 31912 26166 32018 26182
tri 31790 26124 31832 26166 ne
rect 31832 26124 32018 26166
tri 32018 26124 32076 26182 sw
rect 70813 26124 71000 26182
tri 31832 26080 31876 26124 ne
rect 31876 26080 32076 26124
tri 32076 26080 32120 26124 sw
tri 31876 26034 31922 26080 ne
rect 31922 26034 31998 26080
rect 32044 26078 32120 26080
tri 32120 26078 32122 26080 sw
rect 70813 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26034 32122 26078
tri 31922 26020 31936 26034 ne
rect 31936 26020 32122 26034
tri 32122 26020 32180 26078 sw
rect 70813 26020 71000 26078
tri 31936 25974 31982 26020 ne
rect 31982 25974 32180 26020
tri 32180 25974 32226 26020 sw
rect 70813 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
tri 31982 25948 32008 25974 ne
rect 32008 25948 32226 25974
tri 32226 25948 32252 25974 sw
tri 32008 25902 32054 25948 ne
rect 32054 25902 32130 25948
rect 32176 25916 32252 25948
tri 32252 25916 32284 25948 sw
rect 70813 25916 71000 25974
rect 32176 25902 32284 25916
tri 32284 25902 32298 25916 sw
tri 32054 25870 32086 25902 ne
rect 32086 25870 32298 25902
tri 32298 25870 32330 25902 sw
rect 70813 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32086 25816 32140 25870 ne
rect 32140 25816 32330 25870
tri 32140 25770 32186 25816 ne
rect 32186 25770 32262 25816
rect 32308 25812 32330 25816
tri 32330 25812 32388 25870 sw
rect 70813 25812 71000 25870
rect 32308 25770 32388 25812
tri 32186 25766 32190 25770 ne
rect 32190 25766 32388 25770
tri 32388 25766 32434 25812 sw
rect 70813 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
tri 32190 25708 32248 25766 ne
rect 32248 25708 32434 25766
tri 32434 25708 32492 25766 sw
rect 70813 25708 71000 25766
tri 32248 25684 32272 25708 ne
rect 32272 25684 32492 25708
tri 32492 25684 32516 25708 sw
tri 32272 25638 32318 25684 ne
rect 32318 25638 32394 25684
rect 32440 25662 32516 25684
tri 32516 25662 32538 25684 sw
rect 70813 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25638 32538 25662
tri 32318 25604 32352 25638 ne
rect 32352 25604 32538 25638
tri 32538 25604 32596 25662 sw
rect 70813 25604 71000 25662
tri 32352 25558 32398 25604 ne
rect 32398 25558 32596 25604
tri 32596 25558 32642 25604 sw
rect 70813 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
tri 32398 25552 32404 25558 ne
rect 32404 25552 32642 25558
tri 32642 25552 32648 25558 sw
tri 32404 25506 32450 25552 ne
rect 32450 25506 32526 25552
rect 32572 25506 32648 25552
tri 32648 25506 32694 25552 sw
tri 32450 25500 32456 25506 ne
rect 32456 25500 32694 25506
tri 32694 25500 32700 25506 sw
rect 70813 25500 71000 25558
tri 32456 25454 32502 25500 ne
rect 32502 25454 32700 25500
tri 32700 25454 32746 25500 sw
rect 70813 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
tri 32502 25420 32536 25454 ne
rect 32536 25420 32746 25454
tri 32746 25420 32780 25454 sw
tri 32536 25374 32582 25420 ne
rect 32582 25374 32658 25420
rect 32704 25396 32780 25420
tri 32780 25396 32804 25420 sw
rect 70813 25396 71000 25454
rect 32704 25374 32804 25396
tri 32582 25350 32606 25374 ne
rect 32606 25350 32804 25374
tri 32804 25350 32850 25396 sw
rect 70813 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
tri 32606 25292 32664 25350 ne
rect 32664 25292 32850 25350
tri 32850 25292 32908 25350 sw
rect 70813 25292 71000 25350
tri 32664 25288 32668 25292 ne
rect 32668 25288 32908 25292
tri 32908 25288 32912 25292 sw
tri 32668 25242 32714 25288 ne
rect 32714 25242 32790 25288
rect 32836 25246 32912 25288
tri 32912 25246 32954 25288 sw
rect 70813 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 32836 25242 32954 25246
tri 32954 25242 32958 25246 sw
tri 32714 25188 32768 25242 ne
rect 32768 25188 32958 25242
tri 32958 25188 33012 25242 sw
rect 70813 25188 71000 25246
tri 32768 25156 32800 25188 ne
rect 32800 25156 33012 25188
tri 32800 25110 32846 25156 ne
rect 32846 25110 32922 25156
rect 32968 25142 33012 25156
tri 33012 25142 33058 25188 sw
rect 70813 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 32968 25110 33058 25142
tri 32846 25084 32872 25110 ne
rect 32872 25084 33058 25110
tri 33058 25084 33116 25142 sw
rect 70813 25084 71000 25142
tri 32872 25038 32918 25084 ne
rect 32918 25038 33116 25084
tri 33116 25038 33162 25084 sw
rect 70813 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
tri 32918 25024 32932 25038 ne
rect 32932 25024 33162 25038
tri 33162 25024 33176 25038 sw
tri 32932 24978 32978 25024 ne
rect 32978 24978 33054 25024
rect 33100 24980 33176 25024
tri 33176 24980 33220 25024 sw
rect 70813 24980 71000 25038
rect 33100 24978 33220 24980
tri 32978 24934 33022 24978 ne
rect 33022 24934 33220 24978
tri 33220 24934 33266 24980 sw
rect 70813 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33022 24892 33064 24934 ne
rect 33064 24892 33266 24934
tri 33266 24892 33308 24934 sw
tri 33064 24846 33110 24892 ne
rect 33110 24846 33186 24892
rect 33232 24876 33308 24892
tri 33308 24876 33324 24892 sw
rect 70813 24876 71000 24934
rect 33232 24846 33324 24876
tri 33324 24846 33354 24876 sw
tri 33110 24830 33126 24846 ne
rect 33126 24830 33354 24846
tri 33354 24830 33370 24846 sw
rect 70813 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
tri 33126 24772 33184 24830 ne
rect 33184 24772 33370 24830
tri 33370 24772 33428 24830 sw
rect 70813 24772 71000 24830
tri 33184 24760 33196 24772 ne
rect 33196 24760 33428 24772
tri 33196 24714 33242 24760 ne
rect 33242 24714 33318 24760
rect 33364 24726 33428 24760
tri 33428 24726 33474 24772 sw
rect 70813 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 33364 24714 33474 24726
tri 33242 24668 33288 24714 ne
rect 33288 24668 33474 24714
tri 33474 24668 33532 24726 sw
rect 70813 24668 71000 24726
tri 33288 24628 33328 24668 ne
rect 33328 24628 33532 24668
tri 33532 24628 33572 24668 sw
tri 33328 24582 33374 24628 ne
rect 33374 24582 33450 24628
rect 33496 24622 33572 24628
tri 33572 24622 33578 24628 sw
rect 70813 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24582 33578 24622
tri 33578 24582 33618 24622 sw
tri 33374 24564 33392 24582 ne
rect 33392 24564 33618 24582
tri 33618 24564 33636 24582 sw
rect 70813 24564 71000 24622
tri 33392 24518 33438 24564 ne
rect 33438 24518 33636 24564
tri 33636 24518 33682 24564 sw
rect 70813 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33438 24496 33460 24518 ne
rect 33460 24496 33682 24518
tri 33460 24450 33506 24496 ne
rect 33506 24450 33582 24496
rect 33628 24460 33682 24496
tri 33682 24460 33740 24518 sw
rect 70813 24460 71000 24518
rect 33628 24450 33740 24460
tri 33506 24414 33542 24450 ne
rect 33542 24414 33740 24450
tri 33740 24414 33786 24460 sw
rect 70813 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33542 24364 33592 24414 ne
rect 33592 24364 33786 24414
tri 33786 24364 33836 24414 sw
tri 33592 24318 33638 24364 ne
rect 33638 24318 33714 24364
rect 33760 24356 33836 24364
tri 33836 24356 33844 24364 sw
rect 70813 24356 71000 24414
rect 33760 24318 33844 24356
tri 33638 24310 33646 24318 ne
rect 33646 24310 33844 24318
tri 33844 24310 33890 24356 sw
rect 70813 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
tri 33646 24252 33704 24310 ne
rect 33704 24252 33890 24310
tri 33890 24252 33948 24310 sw
rect 70813 24252 71000 24310
tri 33704 24232 33724 24252 ne
rect 33724 24232 33948 24252
tri 33948 24232 33968 24252 sw
tri 33724 24186 33770 24232 ne
rect 33770 24186 33846 24232
rect 33892 24206 33968 24232
tri 33968 24206 33994 24232 sw
rect 70813 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 33892 24186 33994 24206
tri 33994 24186 34014 24206 sw
tri 33770 24148 33808 24186 ne
rect 33808 24148 34014 24186
tri 34014 24148 34052 24186 sw
rect 70813 24148 71000 24206
tri 33808 24102 33854 24148 ne
rect 33854 24102 34052 24148
tri 34052 24102 34098 24148 sw
rect 70813 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
tri 33854 24100 33856 24102 ne
rect 33856 24100 34098 24102
tri 33856 24054 33902 24100 ne
rect 33902 24054 33978 24100
rect 34024 24054 34098 24100
tri 33902 24044 33912 24054 ne
rect 33912 24044 34098 24054
tri 34098 24044 34156 24102 sw
rect 70813 24044 71000 24102
tri 33912 23998 33958 24044 ne
rect 33958 23998 34156 24044
tri 34156 23998 34202 24044 sw
rect 70813 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33958 23968 33988 23998 ne
rect 33988 23968 34202 23998
tri 34202 23968 34232 23998 sw
tri 33988 23922 34034 23968 ne
rect 34034 23922 34110 23968
rect 34156 23940 34232 23968
tri 34232 23940 34260 23968 sw
rect 70813 23940 71000 23998
rect 34156 23922 34260 23940
tri 34034 23894 34062 23922 ne
rect 34062 23894 34260 23922
tri 34260 23894 34306 23940 sw
rect 70813 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34062 23836 34120 23894 ne
rect 34120 23836 34306 23894
tri 34306 23836 34364 23894 sw
rect 70813 23836 71000 23894
tri 34120 23790 34166 23836 ne
rect 34166 23790 34242 23836
rect 34288 23790 34364 23836
tri 34364 23790 34410 23836 sw
rect 70813 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
tri 34166 23732 34224 23790 ne
rect 34224 23732 34410 23790
tri 34410 23732 34468 23790 sw
rect 70813 23732 71000 23790
tri 34224 23704 34252 23732 ne
rect 34252 23704 34468 23732
tri 34468 23704 34496 23732 sw
tri 34252 23658 34298 23704 ne
rect 34298 23658 34374 23704
rect 34420 23686 34496 23704
tri 34496 23686 34514 23704 sw
rect 70813 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23658 34514 23686
tri 34298 23628 34328 23658 ne
rect 34328 23628 34514 23658
tri 34514 23628 34572 23686 sw
rect 70813 23628 71000 23686
tri 34328 23582 34374 23628 ne
rect 34374 23582 34572 23628
tri 34572 23582 34618 23628 sw
rect 70813 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
tri 34374 23572 34384 23582 ne
rect 34384 23572 34618 23582
tri 34618 23572 34628 23582 sw
tri 34384 23526 34430 23572 ne
rect 34430 23526 34506 23572
rect 34552 23526 34628 23572
tri 34628 23526 34674 23572 sw
tri 34430 23524 34432 23526 ne
rect 34432 23524 34674 23526
tri 34674 23524 34676 23526 sw
rect 70813 23524 71000 23582
tri 34432 23478 34478 23524 ne
rect 34478 23478 34676 23524
tri 34676 23478 34722 23524 sw
rect 70813 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
tri 34478 23440 34516 23478 ne
rect 34516 23440 34722 23478
tri 34516 23394 34562 23440 ne
rect 34562 23394 34638 23440
rect 34684 23420 34722 23440
tri 34722 23420 34780 23478 sw
rect 70813 23420 71000 23478
rect 34684 23394 34780 23420
tri 34562 23374 34582 23394 ne
rect 34582 23374 34780 23394
tri 34780 23374 34826 23420 sw
rect 70813 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34582 23316 34640 23374 ne
rect 34640 23316 34826 23374
tri 34826 23316 34884 23374 sw
rect 70813 23316 71000 23374
tri 34640 23308 34648 23316 ne
rect 34648 23308 34884 23316
tri 34884 23308 34892 23316 sw
tri 34648 23262 34694 23308 ne
rect 34694 23262 34770 23308
rect 34816 23270 34892 23308
tri 34892 23270 34930 23308 sw
rect 70813 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 34816 23262 34930 23270
tri 34694 23212 34744 23262 ne
rect 34744 23212 34930 23262
tri 34930 23212 34988 23270 sw
rect 70813 23212 71000 23270
tri 34744 23176 34780 23212 ne
rect 34780 23176 34988 23212
tri 34988 23176 35024 23212 sw
tri 34780 23130 34826 23176 ne
rect 34826 23130 34902 23176
rect 34948 23166 35024 23176
tri 35024 23166 35034 23176 sw
rect 70813 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 34948 23130 35034 23166
tri 35034 23130 35070 23166 sw
tri 34826 23108 34848 23130 ne
rect 34848 23108 35070 23130
tri 35070 23108 35092 23130 sw
rect 70813 23108 71000 23166
tri 34848 23062 34894 23108 ne
rect 34894 23062 35092 23108
tri 35092 23062 35138 23108 sw
rect 70813 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
tri 34894 23044 34912 23062 ne
rect 34912 23044 35138 23062
tri 34912 22998 34958 23044 ne
rect 34958 22998 35034 23044
rect 35080 23004 35138 23044
tri 35138 23004 35196 23062 sw
rect 70813 23004 71000 23062
rect 35080 22998 35196 23004
tri 34958 22958 34998 22998 ne
rect 34998 22958 35196 22998
tri 35196 22958 35242 23004 sw
rect 70813 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 34998 22912 35044 22958 ne
rect 35044 22912 35242 22958
tri 35242 22912 35288 22958 sw
tri 35044 22866 35090 22912 ne
rect 35090 22866 35166 22912
rect 35212 22900 35288 22912
tri 35288 22900 35300 22912 sw
rect 70813 22900 71000 22958
rect 35212 22866 35300 22900
tri 35300 22866 35334 22900 sw
tri 35090 22854 35102 22866 ne
rect 35102 22854 35334 22866
tri 35334 22854 35346 22866 sw
rect 70813 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
tri 35102 22796 35160 22854 ne
rect 35160 22796 35346 22854
tri 35346 22796 35404 22854 sw
rect 70813 22796 71000 22854
tri 35160 22780 35176 22796 ne
rect 35176 22780 35404 22796
tri 35176 22734 35222 22780 ne
rect 35222 22734 35298 22780
rect 35344 22750 35404 22780
tri 35404 22750 35450 22796 sw
rect 70813 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 35344 22734 35450 22750
tri 35222 22692 35264 22734 ne
rect 35264 22692 35450 22734
tri 35450 22692 35508 22750 sw
rect 70813 22692 71000 22750
tri 35264 22648 35308 22692 ne
rect 35308 22648 35508 22692
tri 35508 22648 35552 22692 sw
tri 35308 22602 35354 22648 ne
rect 35354 22602 35430 22648
rect 35476 22646 35552 22648
tri 35552 22646 35554 22648 sw
rect 70813 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22602 35554 22646
tri 35354 22588 35368 22602 ne
rect 35368 22588 35554 22602
tri 35554 22588 35612 22646 sw
rect 70813 22588 71000 22646
tri 35368 22542 35414 22588 ne
rect 35414 22542 35612 22588
tri 35612 22542 35658 22588 sw
rect 70813 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35414 22516 35440 22542 ne
rect 35440 22516 35658 22542
tri 35658 22516 35684 22542 sw
tri 35440 22470 35486 22516 ne
rect 35486 22470 35562 22516
rect 35608 22484 35684 22516
tri 35684 22484 35716 22516 sw
rect 70813 22484 71000 22542
rect 35608 22470 35716 22484
tri 35716 22470 35730 22484 sw
tri 35486 22438 35518 22470 ne
rect 35518 22438 35730 22470
tri 35730 22438 35762 22470 sw
rect 70813 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35518 22384 35572 22438 ne
rect 35572 22384 35762 22438
tri 35572 22338 35618 22384 ne
rect 35618 22338 35694 22384
rect 35740 22380 35762 22384
tri 35762 22380 35820 22438 sw
rect 70813 22380 71000 22438
rect 35740 22338 35820 22380
tri 35618 22334 35622 22338 ne
rect 35622 22334 35820 22338
tri 35820 22334 35866 22380 sw
rect 70813 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35622 22276 35680 22334 ne
rect 35680 22276 35866 22334
tri 35866 22276 35924 22334 sw
rect 70813 22276 71000 22334
tri 35680 22252 35704 22276 ne
rect 35704 22252 35924 22276
tri 35924 22252 35948 22276 sw
tri 35704 22206 35750 22252 ne
rect 35750 22206 35826 22252
rect 35872 22230 35948 22252
tri 35948 22230 35970 22252 sw
rect 70813 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22206 35970 22230
tri 35750 22172 35784 22206 ne
rect 35784 22172 35970 22206
tri 35970 22172 36028 22230 sw
rect 70813 22172 71000 22230
tri 35784 22126 35830 22172 ne
rect 35830 22126 36028 22172
tri 36028 22126 36074 22172 sw
rect 70813 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
tri 35830 22120 35836 22126 ne
rect 35836 22120 36074 22126
tri 36074 22120 36080 22126 sw
tri 35836 22074 35882 22120 ne
rect 35882 22074 35958 22120
rect 36004 22074 36080 22120
tri 36080 22074 36126 22120 sw
tri 35882 22068 35888 22074 ne
rect 35888 22068 36126 22074
tri 36126 22068 36132 22074 sw
rect 70813 22068 71000 22126
tri 35888 22022 35934 22068 ne
rect 35934 22022 36132 22068
tri 36132 22022 36178 22068 sw
rect 70813 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35934 21988 35968 22022 ne
rect 35968 21988 36178 22022
tri 36178 21988 36212 22022 sw
tri 35968 21942 36014 21988 ne
rect 36014 21942 36090 21988
rect 36136 21964 36212 21988
tri 36212 21964 36236 21988 sw
rect 70813 21964 71000 22022
rect 36136 21942 36236 21964
tri 36014 21918 36038 21942 ne
rect 36038 21918 36236 21942
tri 36236 21918 36282 21964 sw
rect 70813 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
tri 36038 21860 36096 21918 ne
rect 36096 21860 36282 21918
tri 36282 21860 36340 21918 sw
rect 70813 21860 71000 21918
tri 36096 21856 36100 21860 ne
rect 36100 21856 36340 21860
tri 36340 21856 36344 21860 sw
tri 36100 21810 36146 21856 ne
rect 36146 21810 36222 21856
rect 36268 21814 36344 21856
tri 36344 21814 36386 21856 sw
rect 70813 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 36268 21810 36386 21814
tri 36386 21810 36390 21814 sw
tri 36146 21756 36200 21810 ne
rect 36200 21756 36390 21810
tri 36390 21756 36444 21810 sw
rect 70813 21756 71000 21814
tri 36200 21724 36232 21756 ne
rect 36232 21724 36444 21756
tri 36232 21678 36278 21724 ne
rect 36278 21678 36354 21724
rect 36400 21710 36444 21724
tri 36444 21710 36490 21756 sw
rect 70813 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 36400 21678 36490 21710
tri 36278 21652 36304 21678 ne
rect 36304 21652 36490 21678
tri 36490 21652 36548 21710 sw
rect 70813 21652 71000 21710
tri 36304 21606 36350 21652 ne
rect 36350 21606 36548 21652
tri 36548 21606 36594 21652 sw
rect 70813 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
tri 36350 21592 36364 21606 ne
rect 36364 21592 36594 21606
tri 36594 21592 36608 21606 sw
tri 36364 21546 36410 21592 ne
rect 36410 21546 36486 21592
rect 36532 21548 36608 21592
tri 36608 21548 36652 21592 sw
rect 70813 21548 71000 21606
rect 36532 21546 36652 21548
tri 36410 21502 36454 21546 ne
rect 36454 21502 36652 21546
tri 36652 21502 36698 21548 sw
rect 70813 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36454 21460 36496 21502 ne
rect 36496 21460 36698 21502
tri 36698 21460 36740 21502 sw
tri 36496 21414 36542 21460 ne
rect 36542 21414 36618 21460
rect 36664 21444 36740 21460
tri 36740 21444 36756 21460 sw
rect 70813 21444 71000 21502
rect 36664 21414 36756 21444
tri 36756 21414 36786 21444 sw
tri 36542 21398 36558 21414 ne
rect 36558 21398 36786 21414
tri 36786 21398 36802 21414 sw
rect 70813 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36558 21340 36616 21398 ne
rect 36616 21340 36802 21398
tri 36802 21340 36860 21398 sw
rect 70813 21340 71000 21398
tri 36616 21328 36628 21340 ne
rect 36628 21328 36860 21340
tri 36628 21282 36674 21328 ne
rect 36674 21282 36750 21328
rect 36796 21294 36860 21328
tri 36860 21294 36906 21340 sw
rect 70813 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36796 21282 36906 21294
tri 36674 21236 36720 21282 ne
rect 36720 21236 36906 21282
tri 36906 21236 36964 21294 sw
rect 70813 21236 71000 21294
tri 36720 21196 36760 21236 ne
rect 36760 21196 36964 21236
tri 36964 21196 37004 21236 sw
tri 36760 21150 36806 21196 ne
rect 36806 21150 36882 21196
rect 36928 21190 37004 21196
tri 37004 21190 37010 21196 sw
rect 70813 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21150 37010 21190
tri 37010 21150 37050 21190 sw
tri 36806 21132 36824 21150 ne
rect 36824 21132 37050 21150
tri 37050 21132 37068 21150 sw
rect 70813 21132 71000 21190
tri 36824 21086 36870 21132 ne
rect 36870 21086 37068 21132
tri 37068 21086 37114 21132 sw
rect 70813 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
tri 36870 21064 36892 21086 ne
rect 36892 21064 37114 21086
tri 36892 21018 36938 21064 ne
rect 36938 21018 37014 21064
rect 37060 21028 37114 21064
tri 37114 21028 37172 21086 sw
rect 70813 21028 71000 21086
rect 37060 21018 37172 21028
tri 36938 20982 36974 21018 ne
rect 36974 20982 37172 21018
tri 37172 20982 37218 21028 sw
rect 70813 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 36974 20932 37024 20982 ne
rect 37024 20932 37218 20982
tri 37218 20932 37268 20982 sw
tri 37024 20886 37070 20932 ne
rect 37070 20886 37146 20932
rect 37192 20924 37268 20932
tri 37268 20924 37276 20932 sw
rect 70813 20924 71000 20982
rect 37192 20886 37276 20924
tri 37070 20878 37078 20886 ne
rect 37078 20878 37276 20886
tri 37276 20878 37322 20924 sw
rect 70813 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
tri 37078 20820 37136 20878 ne
rect 37136 20820 37322 20878
tri 37322 20820 37380 20878 sw
rect 70813 20820 71000 20878
tri 37136 20800 37156 20820 ne
rect 37156 20800 37380 20820
tri 37380 20800 37400 20820 sw
tri 37156 20754 37202 20800 ne
rect 37202 20754 37278 20800
rect 37324 20774 37400 20800
tri 37400 20774 37426 20800 sw
rect 70813 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 37324 20754 37426 20774
tri 37426 20754 37446 20774 sw
tri 37202 20716 37240 20754 ne
rect 37240 20716 37446 20754
tri 37446 20716 37484 20754 sw
rect 70813 20716 71000 20774
tri 37240 20670 37286 20716 ne
rect 37286 20670 37484 20716
tri 37484 20670 37530 20716 sw
rect 70813 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
tri 37286 20668 37288 20670 ne
rect 37288 20668 37530 20670
tri 37288 20622 37334 20668 ne
rect 37334 20622 37410 20668
rect 37456 20622 37530 20668
tri 37334 20612 37344 20622 ne
rect 37344 20612 37530 20622
tri 37530 20612 37588 20670 sw
rect 70813 20612 71000 20670
tri 37344 20566 37390 20612 ne
rect 37390 20566 37588 20612
tri 37588 20566 37634 20612 sw
rect 70813 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
tri 37390 20536 37420 20566 ne
rect 37420 20536 37634 20566
tri 37634 20536 37664 20566 sw
tri 37420 20490 37466 20536 ne
rect 37466 20490 37542 20536
rect 37588 20508 37664 20536
tri 37664 20508 37692 20536 sw
rect 70813 20508 71000 20566
rect 37588 20490 37692 20508
tri 37466 20462 37494 20490 ne
rect 37494 20462 37692 20490
tri 37692 20462 37738 20508 sw
rect 70813 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
tri 37494 20404 37552 20462 ne
rect 37552 20404 37738 20462
tri 37738 20404 37796 20462 sw
rect 70813 20404 71000 20462
tri 37552 20358 37598 20404 ne
rect 37598 20358 37674 20404
rect 37720 20358 37796 20404
tri 37796 20358 37842 20404 sw
rect 70813 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37598 20300 37656 20358 ne
rect 37656 20300 37842 20358
tri 37842 20300 37900 20358 sw
rect 70813 20300 71000 20358
tri 37656 20272 37684 20300 ne
rect 37684 20272 37900 20300
tri 37900 20272 37928 20300 sw
tri 37684 20226 37730 20272 ne
rect 37730 20226 37806 20272
rect 37852 20254 37928 20272
tri 37928 20254 37946 20272 sw
rect 70813 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20226 37946 20254
tri 37730 20196 37760 20226 ne
rect 37760 20196 37946 20226
tri 37946 20196 38004 20254 sw
rect 70813 20196 71000 20254
tri 37760 20150 37806 20196 ne
rect 37806 20150 38004 20196
tri 38004 20150 38050 20196 sw
rect 70813 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
tri 37806 20140 37816 20150 ne
rect 37816 20140 38050 20150
tri 38050 20140 38060 20150 sw
tri 37816 20094 37862 20140 ne
rect 37862 20094 37938 20140
rect 37984 20094 38060 20140
tri 38060 20094 38106 20140 sw
tri 37862 20092 37864 20094 ne
rect 37864 20092 38106 20094
tri 38106 20092 38108 20094 sw
rect 70813 20092 71000 20150
tri 37864 20046 37910 20092 ne
rect 37910 20046 38108 20092
tri 38108 20046 38154 20092 sw
rect 70813 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37910 20008 37948 20046 ne
rect 37948 20008 38154 20046
tri 37948 19962 37994 20008 ne
rect 37994 19962 38070 20008
rect 38116 19988 38154 20008
tri 38154 19988 38212 20046 sw
rect 70813 19988 71000 20046
rect 38116 19962 38212 19988
tri 37994 19942 38014 19962 ne
rect 38014 19942 38212 19962
tri 38212 19942 38258 19988 sw
rect 70813 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
tri 38014 19884 38072 19942 ne
rect 38072 19884 38258 19942
tri 38258 19884 38316 19942 sw
rect 70813 19884 71000 19942
tri 38072 19876 38080 19884 ne
rect 38080 19876 38316 19884
tri 38316 19876 38324 19884 sw
tri 38080 19830 38126 19876 ne
rect 38126 19830 38202 19876
rect 38248 19838 38324 19876
tri 38324 19838 38362 19876 sw
rect 70813 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 38248 19830 38362 19838
tri 38126 19780 38176 19830 ne
rect 38176 19780 38362 19830
tri 38362 19780 38420 19838 sw
rect 70813 19780 71000 19838
tri 38176 19744 38212 19780 ne
rect 38212 19744 38420 19780
tri 38420 19744 38456 19780 sw
tri 38212 19698 38258 19744 ne
rect 38258 19698 38334 19744
rect 38380 19734 38456 19744
tri 38456 19734 38466 19744 sw
rect 70813 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 38380 19698 38466 19734
tri 38466 19698 38502 19734 sw
tri 38258 19676 38280 19698 ne
rect 38280 19676 38502 19698
tri 38502 19676 38524 19698 sw
rect 70813 19676 71000 19734
tri 38280 19630 38326 19676 ne
rect 38326 19630 38524 19676
tri 38524 19630 38570 19676 sw
rect 70813 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
tri 38326 19612 38344 19630 ne
rect 38344 19612 38570 19630
tri 38570 19612 38588 19630 sw
tri 38344 19566 38390 19612 ne
rect 38390 19566 38466 19612
rect 38512 19572 38588 19612
tri 38588 19572 38628 19612 sw
rect 70813 19572 71000 19630
rect 38512 19566 38628 19572
tri 38390 19526 38430 19566 ne
rect 38430 19526 38628 19566
tri 38628 19526 38674 19572 sw
rect 70813 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38430 19480 38476 19526 ne
rect 38476 19480 38674 19526
tri 38674 19480 38720 19526 sw
tri 38476 19434 38522 19480 ne
rect 38522 19434 38598 19480
rect 38644 19468 38720 19480
tri 38720 19468 38732 19480 sw
rect 70813 19468 71000 19526
rect 38644 19434 38732 19468
tri 38732 19434 38766 19468 sw
tri 38522 19422 38534 19434 ne
rect 38534 19422 38766 19434
tri 38766 19422 38778 19434 sw
rect 70813 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
tri 38534 19364 38592 19422 ne
rect 38592 19364 38778 19422
tri 38778 19364 38836 19422 sw
rect 70813 19364 71000 19422
tri 38592 19348 38608 19364 ne
rect 38608 19348 38836 19364
tri 38608 19302 38654 19348 ne
rect 38654 19302 38730 19348
rect 38776 19318 38836 19348
tri 38836 19318 38882 19364 sw
rect 70813 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 38776 19302 38882 19318
tri 38654 19260 38696 19302 ne
rect 38696 19260 38882 19302
tri 38882 19260 38940 19318 sw
rect 70813 19260 71000 19318
tri 38696 19216 38740 19260 ne
rect 38740 19216 38940 19260
tri 38940 19216 38984 19260 sw
tri 38740 19170 38786 19216 ne
rect 38786 19170 38862 19216
rect 38908 19214 38984 19216
tri 38984 19214 38986 19216 sw
rect 70813 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19170 38986 19214
tri 38786 19156 38800 19170 ne
rect 38800 19156 38986 19170
tri 38986 19156 39044 19214 sw
rect 70813 19156 71000 19214
tri 38800 19110 38846 19156 ne
rect 38846 19110 39044 19156
tri 39044 19110 39090 19156 sw
rect 70813 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
tri 38846 19084 38872 19110 ne
rect 38872 19084 39090 19110
tri 39090 19084 39116 19110 sw
tri 38872 19038 38918 19084 ne
rect 38918 19038 38994 19084
rect 39040 19052 39116 19084
tri 39116 19052 39148 19084 sw
rect 70813 19052 71000 19110
rect 39040 19038 39148 19052
tri 39148 19038 39162 19052 sw
tri 38918 19006 38950 19038 ne
rect 38950 19006 39162 19038
tri 39162 19006 39194 19038 sw
rect 70813 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
tri 38950 18952 39004 19006 ne
rect 39004 18952 39194 19006
tri 39004 18906 39050 18952 ne
rect 39050 18906 39126 18952
rect 39172 18948 39194 18952
tri 39194 18948 39252 19006 sw
rect 70813 18948 71000 19006
rect 39172 18906 39252 18948
tri 39050 18902 39054 18906 ne
rect 39054 18902 39252 18906
tri 39252 18902 39298 18948 sw
rect 70813 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
tri 39054 18844 39112 18902 ne
rect 39112 18844 39298 18902
tri 39298 18844 39356 18902 sw
rect 70813 18844 71000 18902
tri 39112 18820 39136 18844 ne
rect 39136 18820 39356 18844
tri 39356 18820 39380 18844 sw
tri 39136 18774 39182 18820 ne
rect 39182 18774 39258 18820
rect 39304 18798 39380 18820
tri 39380 18798 39402 18820 sw
rect 70813 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18774 39402 18798
tri 39182 18740 39216 18774 ne
rect 39216 18740 39402 18774
tri 39402 18740 39460 18798 sw
rect 70813 18740 71000 18798
tri 39216 18694 39262 18740 ne
rect 39262 18694 39460 18740
tri 39460 18694 39506 18740 sw
rect 70813 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
tri 39262 18688 39268 18694 ne
rect 39268 18688 39506 18694
tri 39506 18688 39512 18694 sw
tri 39268 18642 39314 18688 ne
rect 39314 18642 39390 18688
rect 39436 18642 39512 18688
tri 39512 18642 39558 18688 sw
tri 39314 18636 39320 18642 ne
rect 39320 18636 39558 18642
tri 39558 18636 39564 18642 sw
rect 70813 18636 71000 18694
tri 39320 18590 39366 18636 ne
rect 39366 18590 39564 18636
tri 39564 18590 39610 18636 sw
rect 70813 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
tri 39366 18556 39400 18590 ne
rect 39400 18556 39610 18590
tri 39610 18556 39644 18590 sw
tri 39400 18510 39446 18556 ne
rect 39446 18510 39522 18556
rect 39568 18532 39644 18556
tri 39644 18532 39668 18556 sw
rect 70813 18532 71000 18590
rect 39568 18510 39668 18532
tri 39446 18486 39470 18510 ne
rect 39470 18486 39668 18510
tri 39668 18486 39714 18532 sw
rect 70813 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
tri 39470 18428 39528 18486 ne
rect 39528 18428 39714 18486
tri 39714 18428 39772 18486 sw
rect 70813 18428 71000 18486
tri 39528 18424 39532 18428 ne
rect 39532 18424 39772 18428
tri 39772 18424 39776 18428 sw
tri 39532 18378 39578 18424 ne
rect 39578 18378 39654 18424
rect 39700 18382 39776 18424
tri 39776 18382 39818 18424 sw
rect 70813 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 39700 18378 39818 18382
tri 39818 18378 39822 18382 sw
tri 39578 18324 39632 18378 ne
rect 39632 18324 39822 18378
tri 39822 18324 39876 18378 sw
rect 70813 18324 71000 18382
tri 39632 18292 39664 18324 ne
rect 39664 18292 39876 18324
tri 39664 18246 39710 18292 ne
rect 39710 18246 39786 18292
rect 39832 18278 39876 18292
tri 39876 18278 39922 18324 sw
rect 70813 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 39832 18246 39922 18278
tri 39710 18220 39736 18246 ne
rect 39736 18220 39922 18246
tri 39922 18220 39980 18278 sw
rect 70813 18220 71000 18278
tri 39736 18174 39782 18220 ne
rect 39782 18174 39980 18220
tri 39980 18174 40026 18220 sw
rect 70813 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
tri 39782 18160 39796 18174 ne
rect 39796 18160 40026 18174
tri 40026 18160 40040 18174 sw
tri 39796 18114 39842 18160 ne
rect 39842 18114 39918 18160
rect 39964 18116 40040 18160
tri 40040 18116 40084 18160 sw
rect 70813 18116 71000 18174
rect 39964 18114 40084 18116
tri 39842 18070 39886 18114 ne
rect 39886 18070 40084 18114
tri 40084 18070 40130 18116 sw
rect 70813 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39886 18028 39928 18070 ne
rect 39928 18028 40130 18070
tri 40130 18028 40172 18070 sw
tri 39928 17982 39974 18028 ne
rect 39974 17982 40050 18028
rect 40096 18012 40172 18028
tri 40172 18012 40188 18028 sw
rect 70813 18012 71000 18070
rect 40096 17982 40188 18012
tri 40188 17982 40218 18012 sw
tri 39974 17966 39990 17982 ne
rect 39990 17966 40218 17982
tri 40218 17966 40234 17982 sw
rect 70813 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
tri 39990 17908 40048 17966 ne
rect 40048 17908 40234 17966
tri 40234 17908 40292 17966 sw
rect 70813 17908 71000 17966
tri 40048 17896 40060 17908 ne
rect 40060 17896 40292 17908
tri 40292 17896 40304 17908 sw
tri 40060 17850 40106 17896 ne
rect 40106 17850 40182 17896
rect 40228 17862 40304 17896
tri 40304 17862 40338 17896 sw
rect 70813 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 40228 17850 40338 17862
tri 40106 17804 40152 17850 ne
rect 40152 17804 40338 17850
tri 40338 17804 40396 17862 sw
rect 70813 17804 71000 17862
tri 40152 17764 40192 17804 ne
rect 40192 17764 40396 17804
tri 40396 17764 40436 17804 sw
tri 40192 17718 40238 17764 ne
rect 40238 17718 40314 17764
rect 40360 17758 40436 17764
tri 40436 17758 40442 17764 sw
rect 70813 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17718 40442 17758
tri 40442 17718 40482 17758 sw
tri 40238 17700 40256 17718 ne
rect 40256 17700 40482 17718
tri 40482 17700 40500 17718 sw
rect 70813 17700 71000 17758
tri 40256 17654 40302 17700 ne
rect 40302 17654 40500 17700
tri 40500 17654 40546 17700 sw
rect 70813 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40302 17632 40324 17654 ne
rect 40324 17632 40546 17654
tri 40324 17586 40370 17632 ne
rect 40370 17586 40446 17632
rect 40492 17596 40546 17632
tri 40546 17596 40604 17654 sw
rect 70813 17596 71000 17654
rect 40492 17586 40604 17596
tri 40370 17550 40406 17586 ne
rect 40406 17550 40604 17586
tri 40604 17550 40650 17596 sw
rect 70813 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
tri 40406 17500 40456 17550 ne
rect 40456 17500 40650 17550
tri 40650 17500 40700 17550 sw
tri 40456 17454 40502 17500 ne
rect 40502 17454 40578 17500
rect 40624 17492 40700 17500
tri 40700 17492 40708 17500 sw
rect 70813 17492 71000 17550
rect 40624 17454 40708 17492
tri 40708 17454 40746 17492 sw
tri 40502 17446 40510 17454 ne
rect 40510 17446 40746 17454
tri 40746 17446 40754 17454 sw
rect 70813 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
tri 40510 17388 40568 17446 ne
rect 40568 17388 40754 17446
tri 40754 17388 40812 17446 sw
rect 70813 17388 71000 17446
tri 40568 17368 40588 17388 ne
rect 40588 17368 40812 17388
tri 40812 17368 40832 17388 sw
tri 40588 17322 40634 17368 ne
rect 40634 17322 40710 17368
rect 40756 17342 40832 17368
tri 40832 17342 40858 17368 sw
rect 70813 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17322 40858 17342
tri 40858 17322 40878 17342 sw
tri 40634 17284 40672 17322 ne
rect 40672 17284 40878 17322
tri 40878 17284 40916 17322 sw
rect 70813 17284 71000 17342
tri 40672 17238 40718 17284 ne
rect 40718 17238 40916 17284
tri 40916 17238 40962 17284 sw
rect 70813 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
tri 40718 17236 40720 17238 ne
rect 40720 17236 40962 17238
tri 40720 17190 40766 17236 ne
rect 40766 17190 40842 17236
rect 40888 17190 40962 17236
tri 40766 17180 40776 17190 ne
rect 40776 17180 40962 17190
tri 40962 17180 41020 17238 sw
rect 70813 17180 71000 17238
tri 40776 17134 40822 17180 ne
rect 40822 17134 41020 17180
tri 41020 17134 41066 17180 sw
rect 70813 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40822 17104 40852 17134 ne
rect 40852 17104 41066 17134
tri 41066 17104 41096 17134 sw
tri 40852 17058 40898 17104 ne
rect 40898 17058 40974 17104
rect 41020 17076 41096 17104
tri 41096 17076 41124 17104 sw
rect 70813 17076 71000 17134
rect 41020 17058 41124 17076
tri 41124 17058 41142 17076 sw
tri 40898 17030 40926 17058 ne
rect 40926 17030 41142 17058
tri 41142 17030 41170 17058 sw
rect 70813 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
tri 40926 17012 40944 17030 ne
rect 40944 17012 41170 17030
tri 40944 16972 40984 17012 ne
rect 40984 16972 41170 17012
tri 41170 16972 41228 17030 sw
rect 70813 16972 71000 17030
tri 40984 16926 41030 16972 ne
rect 41030 16926 41106 16972
rect 41152 16926 41228 16972
tri 41228 16926 41274 16972 sw
rect 70813 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41030 16868 41088 16926 ne
rect 41088 16868 41274 16926
tri 41274 16868 41332 16926 sw
rect 70813 16868 71000 16926
tri 41088 16840 41116 16868 ne
rect 41116 16840 41332 16868
tri 41332 16840 41360 16868 sw
tri 41116 16794 41162 16840 ne
rect 41162 16794 41238 16840
rect 41284 16822 41360 16840
tri 41360 16822 41378 16840 sw
rect 70813 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16794 41378 16822
tri 41162 16764 41192 16794 ne
rect 41192 16764 41378 16794
tri 41378 16764 41436 16822 sw
rect 70813 16764 71000 16822
tri 41192 16718 41238 16764 ne
rect 41238 16718 41436 16764
tri 41436 16718 41482 16764 sw
rect 70813 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
tri 41238 16708 41248 16718 ne
rect 41248 16708 41482 16718
tri 41482 16708 41492 16718 sw
tri 41248 16662 41294 16708 ne
rect 41294 16662 41370 16708
rect 41416 16662 41492 16708
tri 41492 16662 41538 16708 sw
tri 41294 16660 41296 16662 ne
rect 41296 16660 41538 16662
tri 41538 16660 41540 16662 sw
rect 70813 16660 71000 16718
tri 41296 16614 41342 16660 ne
rect 41342 16614 41540 16660
tri 41540 16614 41586 16660 sw
rect 70813 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
tri 41342 16576 41380 16614 ne
rect 41380 16576 41586 16614
tri 41380 16530 41426 16576 ne
rect 41426 16530 41502 16576
rect 41548 16556 41586 16576
tri 41586 16556 41644 16614 sw
rect 70813 16556 71000 16614
rect 41548 16530 41644 16556
tri 41426 16510 41446 16530 ne
rect 41446 16510 41644 16530
tri 41644 16510 41690 16556 sw
rect 70813 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41446 16452 41504 16510 ne
rect 41504 16452 41690 16510
tri 41690 16452 41748 16510 sw
rect 70813 16452 71000 16510
tri 41504 16444 41512 16452 ne
rect 41512 16444 41748 16452
tri 41748 16444 41756 16452 sw
tri 41512 16398 41558 16444 ne
rect 41558 16398 41634 16444
rect 41680 16406 41756 16444
tri 41756 16406 41794 16444 sw
rect 70813 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 41680 16398 41794 16406
tri 41558 16348 41608 16398 ne
rect 41608 16348 41794 16398
tri 41794 16348 41852 16406 sw
rect 70813 16348 71000 16406
tri 41608 16312 41644 16348 ne
rect 41644 16312 41852 16348
tri 41852 16312 41888 16348 sw
tri 41644 16266 41690 16312 ne
rect 41690 16266 41766 16312
rect 41812 16302 41888 16312
tri 41888 16302 41898 16312 sw
rect 70813 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16266 41898 16302
tri 41898 16266 41934 16302 sw
tri 41690 16244 41712 16266 ne
rect 41712 16244 41934 16266
tri 41934 16244 41956 16266 sw
rect 70813 16244 71000 16302
tri 41712 16198 41758 16244 ne
rect 41758 16198 41956 16244
tri 41956 16198 42002 16244 sw
rect 70813 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
tri 41758 16180 41776 16198 ne
rect 41776 16180 42002 16198
tri 42002 16180 42020 16198 sw
tri 41776 16134 41822 16180 ne
rect 41822 16134 41898 16180
rect 41944 16140 42020 16180
tri 42020 16140 42060 16180 sw
rect 70813 16140 71000 16198
rect 41944 16134 42060 16140
tri 41822 16094 41862 16134 ne
rect 41862 16094 42060 16134
tri 42060 16094 42106 16140 sw
rect 70813 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41862 16048 41908 16094 ne
rect 41908 16048 42106 16094
tri 42106 16048 42152 16094 sw
tri 41908 16002 41954 16048 ne
rect 41954 16002 42030 16048
rect 42076 16036 42152 16048
tri 42152 16036 42164 16048 sw
rect 70813 16036 71000 16094
rect 42076 16002 42164 16036
tri 42164 16002 42198 16036 sw
tri 41954 15990 41966 16002 ne
rect 41966 15990 42198 16002
tri 42198 15990 42210 16002 sw
rect 70813 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
tri 41966 15932 42024 15990 ne
rect 42024 15932 42210 15990
tri 42210 15932 42268 15990 sw
rect 70813 15932 71000 15990
tri 42024 15916 42040 15932 ne
rect 42040 15916 42268 15932
tri 42040 15870 42086 15916 ne
rect 42086 15870 42162 15916
rect 42208 15886 42268 15916
tri 42268 15886 42314 15932 sw
rect 70813 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 42208 15870 42314 15886
tri 42086 15828 42128 15870 ne
rect 42128 15828 42314 15870
tri 42314 15828 42372 15886 sw
rect 70813 15828 71000 15886
tri 42128 15784 42172 15828 ne
rect 42172 15792 42372 15828
tri 42372 15792 42408 15828 sw
rect 42172 15784 42408 15792
tri 42172 15738 42218 15784 ne
rect 42218 15738 42294 15784
rect 42340 15782 42408 15784
tri 42408 15782 42418 15792 sw
rect 70813 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15738 42418 15782
tri 42218 15724 42232 15738 ne
rect 42232 15724 42418 15738
tri 42418 15724 42476 15782 sw
rect 70813 15724 71000 15782
tri 42232 15678 42278 15724 ne
rect 42278 15678 42476 15724
tri 42476 15678 42522 15724 sw
rect 70813 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
tri 42278 15652 42304 15678 ne
rect 42304 15652 42522 15678
tri 42522 15652 42548 15678 sw
tri 42304 15606 42350 15652 ne
rect 42350 15606 42426 15652
rect 42472 15620 42548 15652
tri 42548 15620 42580 15652 sw
rect 70813 15620 71000 15678
rect 42472 15606 42580 15620
tri 42580 15606 42594 15620 sw
tri 42350 15574 42382 15606 ne
rect 42382 15574 42594 15606
tri 42594 15574 42626 15606 sw
rect 70813 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
tri 42382 15548 42408 15574 ne
rect 42408 15548 42626 15574
tri 42626 15548 42652 15574 sw
tri 42408 15520 42436 15548 ne
rect 42436 15520 42652 15548
tri 42436 15474 42482 15520 ne
rect 42482 15474 42558 15520
rect 42604 15516 42652 15520
tri 42652 15516 42684 15548 sw
rect 70813 15516 71000 15574
rect 42604 15474 42684 15516
tri 42482 15470 42486 15474 ne
rect 42486 15470 42684 15474
tri 42684 15470 42730 15516 sw
rect 70813 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
tri 42486 15412 42544 15470 ne
rect 42544 15412 42730 15470
tri 42730 15412 42788 15470 sw
rect 70813 15412 71000 15470
tri 42544 15388 42568 15412 ne
rect 42568 15388 42788 15412
tri 42788 15388 42812 15412 sw
tri 42568 15342 42614 15388 ne
rect 42614 15342 42690 15388
rect 42736 15366 42812 15388
tri 42812 15366 42834 15388 sw
rect 70813 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15342 42834 15366
tri 42834 15342 42858 15366 sw
tri 42614 15308 42648 15342 ne
rect 42648 15308 42858 15342
tri 42858 15308 42892 15342 sw
rect 70813 15308 71000 15366
tri 42648 15304 42652 15308 ne
rect 42652 15304 42892 15308
tri 42652 15262 42694 15304 ne
rect 42694 15262 42892 15304
tri 42892 15262 42938 15308 sw
rect 70813 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
tri 42694 15256 42700 15262 ne
rect 42700 15256 42938 15262
tri 42700 15210 42746 15256 ne
rect 42746 15210 42822 15256
rect 42868 15210 42938 15256
tri 42746 15204 42752 15210 ne
rect 42752 15204 42938 15210
tri 42938 15204 42996 15262 sw
rect 70813 15204 71000 15262
tri 42752 15158 42798 15204 ne
rect 42798 15158 42996 15204
tri 42996 15158 43042 15204 sw
rect 70813 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42798 15124 42832 15158 ne
rect 42832 15124 43042 15158
tri 43042 15124 43076 15158 sw
tri 42832 15078 42878 15124 ne
rect 42878 15078 42954 15124
rect 43000 15100 43076 15124
tri 43076 15100 43100 15124 sw
rect 70813 15100 71000 15158
rect 43000 15078 43100 15100
tri 42878 15054 42902 15078 ne
rect 42902 15054 43100 15078
tri 43100 15054 43146 15100 sw
rect 70813 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42902 14996 42960 15054 ne
rect 42960 14996 43146 15054
tri 43146 14996 43204 15054 sw
rect 70813 14996 71000 15054
tri 42960 14992 42964 14996 ne
rect 42964 14992 43204 14996
tri 43204 14992 43208 14996 sw
tri 42964 14946 43010 14992 ne
rect 43010 14946 43086 14992
rect 43132 14950 43208 14992
tri 43208 14950 43250 14992 sw
rect 70813 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 43132 14946 43250 14950
tri 43250 14946 43254 14950 sw
tri 43010 14892 43064 14946 ne
rect 43064 14892 43254 14946
tri 43254 14892 43308 14946 sw
rect 70813 14892 71000 14950
tri 43064 14860 43096 14892 ne
rect 43096 14860 43308 14892
tri 43308 14860 43340 14892 sw
tri 43096 14814 43142 14860 ne
rect 43142 14814 43218 14860
rect 43264 14846 43340 14860
tri 43340 14846 43354 14860 sw
rect 70813 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 43264 14814 43354 14846
tri 43142 14788 43168 14814 ne
rect 43168 14788 43354 14814
tri 43354 14788 43412 14846 sw
rect 70813 14788 71000 14846
tri 43168 14742 43214 14788 ne
rect 43214 14742 43412 14788
tri 43412 14742 43458 14788 sw
rect 70813 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
tri 43214 14728 43228 14742 ne
rect 43228 14728 43458 14742
tri 43458 14728 43472 14742 sw
tri 43228 14682 43274 14728 ne
rect 43274 14682 43350 14728
rect 43396 14684 43472 14728
tri 43472 14684 43516 14728 sw
rect 70813 14684 71000 14742
rect 43396 14682 43516 14684
tri 43516 14682 43518 14684 sw
tri 43274 14638 43318 14682 ne
rect 43318 14638 43518 14682
tri 43518 14638 43562 14682 sw
rect 70813 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43318 14596 43360 14638 ne
rect 43360 14596 43562 14638
tri 43360 14550 43406 14596 ne
rect 43406 14550 43482 14596
rect 43528 14580 43562 14596
tri 43562 14580 43620 14638 sw
rect 70813 14580 71000 14638
rect 43528 14550 43620 14580
tri 43406 14534 43422 14550 ne
rect 43422 14534 43620 14550
tri 43620 14534 43666 14580 sw
rect 70813 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
tri 43422 14476 43480 14534 ne
rect 43480 14476 43666 14534
tri 43666 14476 43724 14534 sw
rect 70813 14476 71000 14534
tri 43480 14464 43492 14476 ne
rect 43492 14464 43724 14476
tri 43724 14464 43736 14476 sw
tri 43492 14418 43538 14464 ne
rect 43538 14418 43614 14464
rect 43660 14430 43736 14464
tri 43736 14430 43770 14464 sw
rect 70813 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 43660 14418 43770 14430
tri 43538 14372 43584 14418 ne
rect 43584 14372 43770 14418
tri 43770 14372 43828 14430 sw
rect 70813 14372 71000 14430
tri 43584 14332 43624 14372 ne
rect 43624 14332 43828 14372
tri 43828 14332 43868 14372 sw
tri 43624 14286 43670 14332 ne
rect 43670 14286 43746 14332
rect 43792 14326 43868 14332
tri 43868 14326 43874 14332 sw
rect 70813 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43792 14286 43874 14326
tri 43874 14286 43914 14326 sw
tri 43670 14268 43688 14286 ne
rect 43688 14268 43914 14286
tri 43914 14268 43932 14286 sw
rect 70813 14268 71000 14326
tri 43688 14222 43734 14268 ne
rect 43734 14222 43932 14268
tri 43932 14222 43978 14268 sw
rect 70813 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43734 14200 43756 14222 ne
rect 43756 14200 43978 14222
tri 43978 14200 44000 14222 sw
tri 43756 14154 43802 14200 ne
rect 43802 14154 43878 14200
rect 43924 14164 44000 14200
tri 44000 14164 44036 14200 sw
rect 70813 14164 71000 14222
rect 43924 14154 44036 14164
tri 43802 14118 43838 14154 ne
rect 43838 14118 44036 14154
tri 44036 14118 44082 14164 sw
rect 70813 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
tri 43838 14068 43888 14118 ne
rect 43888 14068 44082 14118
tri 44082 14068 44132 14118 sw
tri 43888 14022 43934 14068 ne
rect 43934 14022 44010 14068
rect 44056 14060 44132 14068
tri 44132 14060 44140 14068 sw
rect 70813 14060 71000 14118
rect 44056 14022 44140 14060
tri 44140 14022 44178 14060 sw
tri 43934 14014 43942 14022 ne
rect 43942 14014 44178 14022
tri 44178 14014 44186 14022 sw
rect 70813 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
tri 43942 13956 44000 14014 ne
rect 44000 13956 44186 14014
tri 44186 13956 44244 14014 sw
rect 70813 13956 71000 14014
tri 44000 13936 44020 13956 ne
rect 44020 13936 44244 13956
tri 44020 13890 44066 13936 ne
rect 44066 13890 44142 13936
rect 44188 13910 44244 13936
tri 44244 13910 44290 13956 sw
rect 70813 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 44188 13890 44290 13910
tri 44066 13852 44104 13890 ne
rect 44104 13852 44290 13890
tri 44290 13852 44348 13910 sw
rect 70813 13852 71000 13910
tri 44104 13806 44150 13852 ne
rect 44150 13806 44348 13852
tri 44348 13806 44394 13852 sw
rect 70813 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
tri 44150 13804 44152 13806 ne
rect 44152 13804 44394 13806
tri 44394 13804 44396 13806 sw
tri 44152 13758 44198 13804 ne
rect 44198 13758 44274 13804
rect 44320 13758 44396 13804
tri 44396 13758 44442 13804 sw
tri 44198 13748 44208 13758 ne
rect 44208 13748 44442 13758
tri 44442 13748 44452 13758 sw
rect 70813 13748 71000 13806
tri 44208 13702 44254 13748 ne
rect 44254 13702 44452 13748
tri 44452 13702 44498 13748 sw
rect 70813 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
tri 44254 13672 44284 13702 ne
rect 44284 13672 44498 13702
tri 44284 13626 44330 13672 ne
rect 44330 13626 44406 13672
rect 44452 13644 44498 13672
tri 44498 13644 44556 13702 sw
rect 70813 13644 71000 13702
rect 44452 13626 44556 13644
tri 44330 13598 44358 13626 ne
rect 44358 13598 44556 13626
tri 44556 13598 44602 13644 sw
rect 70813 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
tri 44358 13540 44416 13598 ne
rect 44416 13540 44602 13598
tri 44602 13540 44660 13598 sw
rect 70813 13540 71000 13598
tri 44416 13494 44462 13540 ne
rect 44462 13494 44538 13540
rect 44584 13494 44660 13540
tri 44660 13494 44706 13540 sw
rect 70813 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
tri 44462 13436 44520 13494 ne
rect 44520 13436 44706 13494
tri 44706 13436 44764 13494 sw
rect 70813 13436 71000 13494
tri 44520 13408 44548 13436 ne
rect 44548 13408 44764 13436
tri 44764 13408 44792 13436 sw
tri 44548 13362 44594 13408 ne
rect 44594 13362 44670 13408
rect 44716 13390 44792 13408
tri 44792 13390 44810 13408 sw
rect 70813 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13362 44810 13390
tri 44594 13352 44604 13362 ne
rect 44604 13352 44810 13362
tri 44604 13269 44687 13352 ne
rect 44687 13280 44810 13352
tri 44810 13280 44920 13390 sw
rect 70813 13280 71000 13390
rect 44687 13269 71000 13280
tri 44687 13256 44700 13269 ne
rect 44700 13256 45088 13269
tri 44700 13210 44746 13256 ne
rect 44746 13210 44850 13256
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
tri 44746 13165 44791 13210 ne
rect 44791 13165 71000 13210
tri 44791 13119 44837 13165 ne
rect 44837 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
tri 44837 13108 44848 13119 ne
rect 44848 13108 71000 13119
<< metal2 >>
rect 70584 68116 70702 68200
rect 70584 66916 70613 68116
rect 70669 66916 70702 68116
rect 70584 60120 70702 66916
rect 70584 58920 70613 60120
rect 70669 58920 70702 60120
rect 70584 56910 70702 58920
rect 70584 55710 70613 56910
rect 70669 55710 70702 56910
rect 70584 55302 70702 55710
rect 70584 54102 70613 55302
rect 70669 54102 70702 55302
rect 70584 53722 70702 54102
rect 70584 52522 70613 53722
rect 70669 52522 70702 53722
rect 70584 45739 70702 52522
rect 70584 42875 70613 45739
rect 70669 42875 70702 45739
rect 70584 42497 70702 42875
rect 70584 41297 70613 42497
rect 70669 41297 70702 42497
rect 70584 39332 70702 41297
rect 70584 36468 70613 39332
rect 70669 36468 70702 39332
rect 70584 36132 70702 36468
rect 70584 33268 70613 36132
rect 70669 33268 70702 36132
rect 70584 32920 70702 33268
rect 70584 30056 70613 32920
rect 70669 30056 70702 32920
rect 70584 29752 70702 30056
rect 70584 26888 70613 29752
rect 70669 26888 70702 29752
rect 70584 24906 70702 26888
rect 70584 23706 70613 24906
rect 70669 23706 70702 24906
rect 70584 23599 70702 23706
<< via2 >>
rect 70613 66916 70669 68116
rect 70613 58920 70669 60120
rect 70613 55710 70669 56910
rect 70613 54102 70669 55302
rect 70613 52522 70669 53722
rect 70613 42875 70669 45739
rect 70613 41297 70669 42497
rect 70613 36468 70669 39332
rect 70613 33268 70669 36132
rect 70613 30056 70669 32920
rect 70613 26888 70669 29752
rect 70613 23706 70669 24906
<< metal3 >>
rect 14000 47112 17000 71000
rect 17200 48448 20200 71000
rect 20400 49774 23400 71000
rect 23600 50451 25000 71000
rect 25200 51220 26600 71000
rect 26800 52454 29800 71000
rect 30000 53792 33000 71000
rect 33200 55124 36200 71000
rect 36400 56465 39400 71000
rect 39600 57138 41000 71000
rect 41200 57723 42600 71000
rect 42800 59150 45800 71000
rect 46000 60510 49000 71000
rect 49200 61175 50600 71000
rect 50800 61839 52200 71000
rect 52400 62507 53800 71000
rect 54000 63173 55400 71000
rect 55600 63836 57000 71000
rect 57200 64499 58600 71000
rect 58800 65166 60200 71000
rect 60400 65831 61800 71000
rect 62000 66494 63400 71000
rect 63600 67166 65000 71000
rect 65200 67829 66600 71000
rect 66800 68476 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68400 68693 68476 68769 ne
rect 68476 68693 71000 68769
tri 68200 68476 68417 68693 sw
tri 68476 68476 68693 68693 ne
rect 68693 68476 71000 68693
rect 66800 68200 68417 68476
tri 68417 68200 68693 68476 sw
tri 68693 68400 68769 68476 ne
rect 68769 68400 71000 68476
rect 66800 68116 71000 68200
rect 66800 68113 70613 68116
tri 66800 68029 66884 68113 ne
rect 66884 68029 70613 68113
tri 66600 67829 66800 68029 sw
tri 66884 67829 67084 68029 ne
rect 67084 67829 70613 68029
rect 65200 67545 66800 67829
tri 66800 67545 67084 67829 sw
tri 67084 67545 67368 67829 ne
rect 67368 67545 70613 67829
rect 65200 67449 67084 67545
tri 65200 67366 65283 67449 ne
rect 65283 67368 67084 67449
tri 67084 67368 67261 67545 sw
tri 67368 67368 67545 67545 ne
rect 67545 67368 70613 67545
rect 65283 67366 67261 67368
tri 65000 67166 65200 67366 sw
tri 65283 67166 65483 67366 ne
rect 65483 67166 67261 67366
rect 63600 66883 65200 67166
tri 65200 66883 65483 67166 sw
tri 65483 66883 65766 67166 ne
rect 65766 67084 67261 67166
tri 67261 67084 67545 67368 sw
tri 67545 67084 67829 67368 ne
rect 67829 67084 70613 67368
rect 65766 66883 67545 67084
rect 63600 66786 65483 66883
tri 63600 66694 63692 66786 ne
rect 63692 66694 65483 66786
tri 63400 66494 63600 66694 sw
tri 63692 66494 63892 66694 ne
rect 63892 66600 65483 66694
tri 65483 66600 65766 66883 sw
tri 65766 66600 66049 66883 ne
rect 66049 66800 67545 66883
tri 67545 66800 67829 67084 sw
tri 67829 66800 68113 67084 ne
rect 68113 66916 70613 67084
rect 70669 66916 71000 68116
rect 68113 66800 71000 66916
rect 66049 66600 67829 66800
tri 67829 66600 68029 66800 sw
rect 63892 66494 65766 66600
rect 62000 66202 63600 66494
tri 63600 66202 63892 66494 sw
tri 63892 66202 64184 66494 ne
rect 64184 66332 65766 66494
tri 65766 66332 66034 66600 sw
tri 66049 66332 66317 66600 ne
rect 66317 66332 71000 66600
rect 64184 66202 66034 66332
rect 62000 66114 63892 66202
tri 62000 66031 62083 66114 ne
rect 62083 66031 63892 66114
tri 61800 65831 62000 66031 sw
tri 62083 65831 62283 66031 ne
rect 62283 65964 63892 66031
tri 63892 65964 64130 66202 sw
tri 64184 65964 64422 66202 ne
rect 64422 66049 66034 66202
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64422 65964 66317 66049
rect 62283 65831 64130 65964
rect 60400 65663 62000 65831
tri 62000 65663 62168 65831 sw
tri 62283 65663 62451 65831 ne
rect 62451 65672 64130 65831
tri 64130 65672 64422 65964 sw
tri 64422 65672 64714 65964 ne
rect 64714 65766 66317 65964
tri 66317 65766 66600 66049 sw
tri 66600 65766 66883 66049 ne
rect 66883 65766 71000 66049
rect 64714 65672 66600 65766
rect 62451 65663 64422 65672
rect 60400 65451 62168 65663
tri 60400 65366 60485 65451 ne
rect 60485 65380 62168 65451
tri 62168 65380 62451 65663 sw
tri 62451 65380 62734 65663 ne
rect 62734 65380 64422 65663
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65483 66600 65672
tri 66600 65483 66883 65766 sw
tri 66883 65483 67166 65766 ne
rect 67166 65483 71000 65766
rect 65006 65380 66883 65483
rect 60485 65366 62451 65380
tri 60200 65166 60400 65366 sw
tri 60485 65166 60685 65366 ne
rect 60685 65166 62451 65366
rect 58800 64881 60400 65166
tri 60400 64881 60685 65166 sw
tri 60685 64881 60970 65166 ne
rect 60970 65097 62451 65166
tri 62451 65097 62734 65380 sw
tri 62734 65097 63017 65380 ne
rect 63017 65292 64714 65380
tri 64714 65292 64802 65380 sw
tri 65006 65292 65094 65380 ne
rect 65094 65292 66883 65380
rect 63017 65097 64802 65292
rect 60970 64997 62734 65097
tri 62734 64997 62834 65097 sw
tri 63017 64997 63117 65097 ne
rect 63117 65000 64802 65097
tri 64802 65000 65094 65292 sw
tri 65094 65000 65386 65292 ne
rect 65386 65200 66883 65292
tri 66883 65200 67166 65483 sw
tri 67166 65200 67449 65483 ne
rect 67449 65200 71000 65483
rect 65386 65000 67166 65200
tri 67166 65000 67366 65200 sw
rect 63117 64997 65094 65000
rect 60970 64881 62834 64997
rect 58800 64786 60685 64881
tri 58800 64699 58887 64786 ne
rect 58887 64730 60685 64786
tri 60685 64730 60836 64881 sw
tri 60970 64730 61121 64881 ne
rect 61121 64730 62834 64881
rect 58887 64699 60836 64730
tri 58600 64499 58800 64699 sw
tri 58887 64499 59087 64699 ne
rect 59087 64499 60836 64699
rect 57200 64447 58800 64499
tri 58800 64447 58852 64499 sw
tri 59087 64447 59139 64499 ne
rect 59139 64447 60836 64499
rect 57200 64160 58852 64447
tri 58852 64160 59139 64447 sw
tri 59139 64160 59426 64447 ne
rect 59426 64445 60836 64447
tri 60836 64445 61121 64730 sw
tri 61121 64445 61406 64730 ne
rect 61406 64714 62834 64730
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61406 64445 63117 64714
rect 59426 64160 61121 64445
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63117 64445
tri 63117 64431 63400 64714 sw
tri 63400 64431 63683 64714 ne
rect 63683 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63683 64431 65386 64708
rect 61691 64160 63400 64431
rect 57200 64119 59139 64160
tri 57200 64036 57283 64119 ne
rect 57283 64036 59139 64119
tri 57000 63836 57200 64036 sw
tri 57283 63836 57483 64036 ne
rect 57483 63873 59139 64036
tri 59139 63873 59426 64160 sw
tri 59426 63873 59713 64160 ne
rect 59713 64065 61406 64160
tri 61406 64065 61501 64160 sw
tri 61691 64065 61786 64160 ne
rect 61786 64148 63400 64160
tri 63400 64148 63683 64431 sw
tri 63683 64148 63966 64431 ne
rect 63966 64416 65386 64431
tri 65386 64416 65678 64708 sw
tri 65678 64416 65970 64708 ne
rect 65970 64416 71000 64708
rect 63966 64184 65678 64416
tri 65678 64184 65910 64416 sw
tri 65970 64184 66202 64416 ne
rect 66202 64184 71000 64416
rect 63966 64148 65910 64184
rect 61786 64065 63683 64148
rect 59713 63873 61501 64065
rect 57483 63836 59426 63873
rect 55600 63553 57200 63836
tri 57200 63553 57483 63836 sw
tri 57483 63553 57766 63836 ne
rect 57766 63673 59426 63836
tri 59426 63673 59626 63873 sw
tri 59713 63673 59913 63873 ne
rect 59913 63780 61501 63873
tri 61501 63780 61786 64065 sw
tri 61786 63780 62071 64065 ne
rect 62071 63966 63683 64065
tri 63683 63966 63865 64148 sw
tri 63966 63966 64148 64148 ne
rect 64148 63966 65910 64148
rect 62071 63780 63865 63966
rect 59913 63673 61786 63780
rect 57766 63553 59626 63673
rect 55600 63506 57483 63553
tri 57483 63506 57530 63553 sw
tri 57766 63506 57813 63553 ne
rect 57813 63506 59626 63553
rect 55600 63456 57530 63506
tri 55600 63373 55683 63456 ne
rect 55683 63373 57530 63456
tri 55400 63173 55600 63373 sw
tri 55683 63173 55883 63373 ne
rect 55883 63223 57530 63373
tri 57530 63223 57813 63506 sw
tri 57813 63223 58096 63506 ne
rect 58096 63386 59626 63506
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63683 63865 63780
tri 63865 63683 64148 63966 sw
tri 64148 63683 64431 63966 ne
rect 64431 63892 65910 63966
tri 65910 63892 66202 64184 sw
tri 66202 63892 66494 64184 ne
rect 66494 63892 71000 64184
rect 64431 63683 66202 63892
rect 62356 63495 64148 63683
rect 60200 63386 62071 63495
rect 58096 63223 59913 63386
rect 55883 63173 57813 63223
rect 54000 62940 55600 63173
tri 55600 62940 55833 63173 sw
tri 55883 62940 56116 63173 ne
rect 56116 62940 57813 63173
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59913 63223
tri 59913 63099 60200 63386 sw
tri 60200 63099 60487 63386 ne
rect 60487 63210 62071 63386
tri 62071 63210 62356 63495 sw
tri 62356 63210 62641 63495 ne
rect 62641 63400 64148 63495
tri 64148 63400 64431 63683 sw
tri 64431 63400 64714 63683 ne
rect 64714 63600 66202 63683
tri 66202 63600 66494 63892 sw
tri 66494 63600 66786 63892 ne
rect 66786 63600 71000 63892
rect 64714 63400 66494 63600
tri 66494 63400 66694 63600 sw
rect 62641 63210 64431 63400
rect 60487 63099 62356 63210
rect 58379 62940 60200 63099
rect 54000 62793 55833 62940
tri 54000 62707 54086 62793 ne
rect 54086 62707 55833 62793
tri 53800 62507 54000 62707 sw
tri 54086 62507 54286 62707 ne
rect 54286 62657 55833 62707
tri 55833 62657 56116 62940 sw
tri 56116 62657 56399 62940 ne
rect 56399 62843 58096 62940
tri 58096 62843 58193 62940 sw
tri 58379 62843 58476 62940 ne
rect 58476 62843 60200 62940
rect 56399 62657 58193 62843
rect 54286 62622 56116 62657
tri 56116 62622 56151 62657 sw
tri 56399 62622 56434 62657 ne
rect 56434 62622 58193 62657
rect 54286 62507 56151 62622
rect 52400 62221 54000 62507
tri 54000 62221 54286 62507 sw
tri 54286 62221 54572 62507 ne
rect 54572 62339 56151 62507
tri 56151 62339 56434 62622 sw
tri 56434 62339 56717 62622 ne
rect 56717 62560 58193 62622
tri 58193 62560 58476 62843 sw
tri 58476 62560 58759 62843 ne
rect 58759 62812 60200 62843
tri 60200 62812 60487 63099 sw
tri 60487 62812 60774 63099 ne
rect 60774 62925 62356 63099
tri 62356 62925 62641 63210 sw
tri 62641 62925 62926 63210 ne
rect 62926 63117 64431 63210
tri 64431 63117 64714 63400 sw
tri 64714 63117 64997 63400 ne
rect 64997 63117 71000 63400
rect 62926 62925 64714 63117
rect 60774 62812 62641 62925
rect 58759 62754 60487 62812
tri 60487 62754 60545 62812 sw
tri 60774 62754 60832 62812 ne
rect 60832 62754 62641 62812
rect 58759 62560 60545 62754
rect 56717 62339 58476 62560
rect 54572 62221 56434 62339
rect 52400 62127 54286 62221
tri 52400 62039 52488 62127 ne
rect 52488 62039 54286 62127
tri 52200 61839 52400 62039 sw
tri 52488 61839 52688 62039 ne
rect 52688 62006 54286 62039
tri 54286 62006 54501 62221 sw
tri 54572 62006 54787 62221 ne
rect 54787 62056 56434 62221
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62467 60545 62560
tri 60545 62467 60832 62754 sw
tri 60832 62467 61119 62754 ne
rect 61119 62750 62641 62754
tri 62641 62750 62816 62925 sw
tri 62926 62750 63101 62925 ne
rect 63101 62834 64714 62925
tri 64714 62834 64997 63117 sw
tri 64997 62834 65280 63117 ne
rect 65280 62834 71000 63117
rect 63101 62750 64997 62834
rect 61119 62467 62816 62750
rect 59042 62277 60832 62467
rect 57000 62056 58759 62277
rect 54787 62006 56717 62056
rect 52688 61839 54501 62006
rect 50800 61720 52400 61839
tri 52400 61720 52519 61839 sw
tri 52688 61720 52807 61839 ne
rect 52807 61720 54501 61839
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56717 62006
tri 56717 61773 57000 62056 sw
tri 57000 61773 57283 62056 ne
rect 57283 61994 58759 62056
tri 58759 61994 59042 62277 sw
tri 59042 61994 59325 62277 ne
rect 59325 62180 60832 62277
tri 60832 62180 61119 62467 sw
tri 61119 62180 61406 62467 ne
rect 61406 62465 62816 62467
tri 62816 62465 63101 62750 sw
tri 63101 62465 63386 62750 ne
rect 63386 62566 64997 62750
tri 64997 62566 65265 62834 sw
tri 65280 62566 65548 62834 ne
rect 65548 62566 71000 62834
rect 63386 62465 65265 62566
rect 61406 62180 63101 62465
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62283 65265 62465
tri 65265 62283 65548 62566 sw
tri 65548 62283 65831 62566 ne
rect 65831 62283 71000 62566
rect 63671 62180 65548 62283
rect 59325 61994 61119 62180
rect 57283 61773 59042 61994
rect 55073 61720 57000 61773
rect 50800 61459 52519 61720
tri 50800 61375 50884 61459 ne
rect 50884 61432 52519 61459
tri 52519 61432 52807 61720 sw
tri 52807 61432 53095 61720 ne
rect 53095 61626 54787 61720
tri 54787 61626 54881 61720 sw
tri 55073 61626 55167 61720 ne
rect 55167 61626 57000 61720
rect 53095 61432 54881 61626
rect 50884 61375 52807 61432
tri 50600 61175 50800 61375 sw
tri 50884 61175 51084 61375 ne
rect 51084 61303 52807 61375
tri 52807 61303 52936 61432 sw
tri 53095 61303 53224 61432 ne
rect 53224 61340 54881 61432
tri 54881 61340 55167 61626 sw
tri 55167 61340 55453 61626 ne
rect 55453 61490 57000 61626
tri 57000 61490 57283 61773 sw
tri 57283 61490 57566 61773 ne
rect 57566 61711 59042 61773
tri 59042 61711 59325 61994 sw
tri 59325 61711 59608 61994 ne
rect 59608 61893 61119 61994
tri 61119 61893 61406 62180 sw
tri 61406 61893 61693 62180 ne
rect 61693 62085 63386 62180
tri 63386 62085 63481 62180 sw
tri 63671 62085 63766 62180 ne
rect 63766 62085 65548 62180
rect 61693 61893 63481 62085
rect 59608 61711 61406 61893
rect 57566 61526 59325 61711
tri 59325 61526 59510 61711 sw
tri 59608 61526 59793 61711 ne
rect 59793 61606 61406 61711
tri 61406 61606 61693 61893 sw
tri 61693 61606 61980 61893 ne
rect 61980 61800 63481 61893
tri 63481 61800 63766 62085 sw
tri 63766 61800 64051 62085 ne
rect 64051 62000 65548 62085
tri 65548 62000 65831 62283 sw
tri 65831 62000 66114 62283 ne
rect 66114 62000 71000 62283
rect 64051 61800 65831 62000
tri 65831 61800 66031 62000 sw
rect 61980 61606 63766 61800
rect 59793 61526 61693 61606
rect 57566 61490 59510 61526
rect 55453 61340 57283 61490
rect 53224 61303 55167 61340
rect 51084 61175 52936 61303
rect 49200 60891 50800 61175
tri 50800 60891 51084 61175 sw
tri 51084 60891 51368 61175 ne
rect 51368 61015 52936 61175
tri 52936 61015 53224 61303 sw
tri 53224 61015 53512 61303 ne
rect 53512 61054 55167 61303
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61243 57283 61340
tri 57283 61243 57530 61490 sw
tri 57566 61243 57813 61490 ne
rect 57813 61243 59510 61490
tri 59510 61243 59793 61526 sw
tri 59793 61243 60076 61526 ne
rect 60076 61319 61693 61526
tri 61693 61319 61980 61606 sw
tri 61980 61319 62267 61606 ne
rect 62267 61515 63766 61606
tri 63766 61515 64051 61800 sw
tri 64051 61515 64336 61800 ne
rect 64336 61515 71000 61800
rect 62267 61319 64051 61515
rect 60076 61243 61980 61319
rect 55739 61054 57530 61243
rect 53512 61015 55453 61054
rect 51368 60891 53224 61015
rect 49200 60795 51084 60891
tri 49200 60710 49285 60795 ne
rect 49285 60784 51084 60795
tri 51084 60784 51191 60891 sw
tri 51368 60784 51475 60891 ne
rect 51475 60784 53224 60891
rect 49285 60710 51191 60784
tri 49000 60510 49200 60710 sw
tri 49285 60510 49485 60710 ne
rect 49485 60510 51191 60710
rect 46000 60500 49200 60510
tri 49200 60500 49210 60510 sw
tri 49485 60500 49495 60510 ne
rect 49495 60500 51191 60510
tri 51191 60500 51475 60784 sw
tri 51475 60500 51759 60784 ne
rect 51759 60727 53224 60784
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60768 55453 61015
tri 55453 60768 55739 61054 sw
tri 55739 60768 56025 61054 ne
rect 56025 60960 57530 61054
tri 57530 60960 57813 61243 sw
tri 57813 60960 58096 61243 ne
rect 58096 60960 59793 61243
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 61154 61980 61243
tri 61980 61154 62145 61319 sw
tri 62267 61154 62432 61319 ne
rect 62432 61230 64051 61319
tri 64051 61230 64336 61515 sw
tri 64336 61230 64621 61515 ne
rect 64621 61230 71000 61515
rect 62432 61154 64336 61230
rect 60359 60960 62145 61154
rect 56025 60768 57813 60960
rect 53800 60727 55739 60768
rect 51759 60500 53512 60727
rect 46000 60215 49210 60500
tri 49210 60215 49495 60500 sw
tri 49495 60215 49780 60500 ne
rect 49780 60404 51475 60500
tri 51475 60404 51571 60500 sw
tri 51759 60404 51855 60500 ne
rect 51855 60439 53512 60500
tri 53512 60439 53800 60727 sw
tri 53800 60439 54088 60727 ne
rect 54088 60482 55739 60727
tri 55739 60482 56025 60768 sw
tri 56025 60482 56311 60768 ne
rect 56311 60677 57813 60768
tri 57813 60677 58096 60960 sw
tri 58096 60677 58379 60960 ne
rect 58379 60863 60076 60960
tri 60076 60863 60173 60960 sw
tri 60359 60863 60456 60960 ne
rect 60456 60867 62145 60960
tri 62145 60867 62432 61154 sw
tri 62432 60867 62719 61154 ne
rect 62719 60970 64336 61154
tri 64336 60970 64596 61230 sw
tri 64621 60970 64881 61230 ne
rect 64881 60970 71000 61230
rect 62719 60867 64596 60970
rect 60456 60863 62432 60867
rect 58379 60677 60173 60863
rect 56311 60482 58096 60677
rect 54088 60439 56025 60482
rect 51855 60404 53800 60439
rect 49780 60215 51571 60404
rect 46000 59965 49495 60215
tri 49495 59965 49745 60215 sw
tri 49780 59965 50030 60215 ne
rect 50030 60120 51571 60215
tri 51571 60120 51855 60404 sw
tri 51855 60120 52139 60404 ne
rect 52139 60151 53800 60404
tri 53800 60151 54088 60439 sw
tri 54088 60151 54376 60439 ne
rect 54376 60312 56025 60439
tri 56025 60312 56195 60482 sw
tri 56311 60312 56481 60482 ne
rect 56481 60394 58096 60482
tri 58096 60394 58379 60677 sw
tri 58379 60394 58662 60677 ne
rect 58662 60580 60173 60677
tri 60173 60580 60456 60863 sw
tri 60456 60580 60739 60863 ne
rect 60739 60580 62432 60863
tri 62432 60580 62719 60867 sw
tri 62719 60580 63006 60867 ne
rect 63006 60685 64596 60867
tri 64596 60685 64881 60970 sw
tri 64881 60685 65166 60970 ne
rect 65166 60685 71000 60970
rect 63006 60580 64881 60685
rect 58662 60394 60456 60580
rect 56481 60312 58379 60394
rect 54376 60151 56195 60312
rect 52139 60120 54088 60151
rect 50030 60059 51855 60120
tri 51855 60059 51916 60120 sw
tri 52139 60059 52200 60120 ne
rect 52200 60059 54088 60120
rect 50030 59965 51916 60059
rect 46000 59680 49745 59965
tri 49745 59680 50030 59965 sw
tri 50030 59680 50315 59965 ne
rect 50315 59775 51916 59965
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 60028 54088 60059
tri 54088 60028 54211 60151 sw
tri 54376 60028 54499 60151 ne
rect 54499 60028 56195 60151
rect 52484 59775 54211 60028
rect 50315 59680 52200 59775
rect 46000 59461 50030 59680
tri 46000 59350 46111 59461 ne
rect 46111 59395 50030 59461
tri 50030 59395 50315 59680 sw
tri 50315 59395 50600 59680 ne
rect 50600 59491 52200 59680
tri 52200 59491 52484 59775 sw
tri 52484 59491 52768 59775 ne
rect 52768 59740 54211 59775
tri 54211 59740 54499 60028 sw
tri 54499 59740 54787 60028 ne
rect 54787 60026 56195 60028
tri 56195 60026 56481 60312 sw
tri 56481 60026 56767 60312 ne
rect 56767 60111 58379 60312
tri 58379 60111 58662 60394 sw
tri 58662 60111 58945 60394 ne
rect 58945 60297 60456 60394
tri 60456 60297 60739 60580 sw
tri 60739 60297 61022 60580 ne
rect 61022 60487 62719 60580
tri 62719 60487 62812 60580 sw
tri 63006 60487 63099 60580 ne
rect 63099 60487 64881 60580
rect 61022 60297 62812 60487
rect 58945 60111 60739 60297
rect 56767 60026 58662 60111
rect 54787 59740 56481 60026
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 59926 58662 60026
tri 58662 59926 58847 60111 sw
tri 58945 59926 59130 60111 ne
rect 59130 60014 60739 60111
tri 60739 60014 61022 60297 sw
tri 61022 60014 61305 60297 ne
rect 61305 60200 62812 60297
tri 62812 60200 63099 60487 sw
tri 63099 60200 63386 60487 ne
rect 63386 60400 64881 60487
tri 64881 60400 65166 60685 sw
tri 65166 60400 65451 60685 ne
rect 65451 60400 71000 60685
rect 63386 60200 65166 60400
tri 65166 60200 65366 60400 sw
rect 61305 60014 63099 60200
rect 59130 59926 61022 60014
rect 57053 59740 58847 59926
rect 52768 59491 54499 59740
rect 50600 59395 52484 59491
rect 46111 59350 50315 59395
tri 45800 59150 46000 59350 sw
tri 46111 59150 46311 59350 ne
rect 46311 59150 50315 59350
rect 42800 58920 46000 59150
tri 46000 58920 46230 59150 sw
tri 46311 58920 46541 59150 ne
rect 46541 59110 50315 59150
tri 50315 59110 50600 59395 sw
tri 50600 59110 50885 59395 ne
rect 50885 59207 52484 59395
tri 52484 59207 52768 59491 sw
tri 52768 59207 53052 59491 ne
rect 53052 59452 54499 59491
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59646 56767 59740
tri 56767 59646 56861 59740 sw
tri 57053 59646 57147 59740 ne
rect 57147 59646 58847 59740
rect 55075 59452 56861 59646
rect 53052 59207 54787 59452
rect 50885 59110 52768 59207
rect 46541 58920 50600 59110
rect 42800 58747 46230 58920
tri 46230 58747 46403 58920 sw
tri 46541 58747 46714 58920 ne
rect 46714 58825 50600 58920
tri 50600 58825 50885 59110 sw
tri 50885 58825 51170 59110 ne
rect 51170 59088 52768 59110
tri 52768 59088 52887 59207 sw
tri 53052 59088 53171 59207 ne
rect 53171 59164 54787 59207
tri 54787 59164 55075 59452 sw
tri 55075 59164 55363 59452 ne
rect 55363 59360 56861 59452
tri 56861 59360 57147 59646 sw
tri 57147 59360 57433 59646 ne
rect 57433 59643 58847 59646
tri 58847 59643 59130 59926 sw
tri 59130 59643 59413 59926 ne
rect 59413 59731 61022 59926
tri 61022 59731 61305 60014 sw
tri 61305 59731 61588 60014 ne
rect 61588 59913 63099 60014
tri 63099 59913 63386 60200 sw
tri 63386 59913 63673 60200 ne
rect 63673 60120 71000 60200
rect 63673 59913 70613 60120
rect 61588 59731 63386 59913
rect 59413 59643 61305 59731
rect 57433 59360 59130 59643
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59546 61305 59643
tri 61305 59546 61490 59731 sw
tri 61588 59546 61773 59731 ne
rect 61773 59626 63386 59731
tri 63386 59626 63673 59913 sw
tri 63673 59626 63960 59913 ne
rect 63960 59626 70613 59913
rect 61773 59546 63673 59626
rect 59696 59360 61490 59546
rect 55363 59164 57147 59360
rect 53171 59088 55075 59164
rect 51170 58825 52887 59088
rect 46714 58805 50885 58825
tri 50885 58805 50905 58825 sw
tri 51170 58805 51190 58825 ne
rect 51190 58805 52887 58825
rect 46714 58747 50905 58805
rect 42800 58436 46403 58747
tri 46403 58436 46714 58747 sw
tri 46714 58436 47025 58747 ne
rect 47025 58520 50905 58747
tri 50905 58520 51190 58805 sw
tri 51190 58520 51475 58805 ne
rect 51475 58804 52887 58805
tri 52887 58804 53171 59088 sw
tri 53171 58804 53455 59088 ne
rect 53455 58876 55075 59088
tri 55075 58876 55363 59164 sw
tri 55363 58876 55651 59164 ne
rect 55651 59074 57147 59164
tri 57147 59074 57433 59360 sw
tri 57433 59074 57719 59360 ne
rect 57719 59263 59413 59360
tri 59413 59263 59510 59360 sw
tri 59696 59263 59793 59360 ne
rect 59793 59263 61490 59360
tri 61490 59263 61773 59546 sw
tri 61773 59263 62056 59546 ne
rect 62056 59374 63673 59546
tri 63673 59374 63925 59626 sw
tri 63960 59374 64212 59626 ne
rect 64212 59374 70613 59626
rect 62056 59263 63925 59374
rect 57719 59074 59510 59263
rect 55651 58876 57433 59074
rect 53455 58804 55363 58876
rect 51475 58520 53171 58804
tri 53171 58520 53455 58804 sw
tri 53455 58520 53739 58804 ne
rect 53739 58716 55363 58804
tri 55363 58716 55523 58876 sw
tri 55651 58716 55811 58876 ne
rect 55811 58788 57433 58876
tri 57433 58788 57719 59074 sw
tri 57719 58788 58005 59074 ne
rect 58005 58980 59510 59074
tri 59510 58980 59793 59263 sw
tri 59793 58980 60076 59263 ne
rect 60076 58980 61773 59263
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 59087 63925 59263
tri 63925 59087 64212 59374 sw
tri 64212 59087 64499 59374 ne
rect 64499 59087 70613 59374
rect 62339 58980 64212 59087
rect 58005 58788 59793 58980
rect 55811 58716 57719 58788
rect 53739 58520 55523 58716
rect 47025 58436 51190 58520
rect 42800 58125 46714 58436
tri 46714 58125 47025 58436 sw
tri 47025 58125 47336 58436 ne
rect 47336 58235 51190 58436
tri 51190 58235 51475 58520 sw
tri 51475 58235 51760 58520 ne
rect 51760 58424 53455 58520
tri 53455 58424 53551 58520 sw
tri 53739 58424 53835 58520 ne
rect 53835 58428 55523 58520
tri 55523 58428 55811 58716 sw
tri 55811 58428 56099 58716 ne
rect 56099 58502 57719 58716
tri 57719 58502 58005 58788 sw
tri 58005 58502 58291 58788 ne
rect 58291 58697 59793 58788
tri 59793 58697 60076 58980 sw
tri 60076 58697 60359 58980 ne
rect 60359 58883 62056 58980
tri 62056 58883 62153 58980 sw
tri 62339 58883 62436 58980 ne
rect 62436 58883 64212 58980
rect 60359 58697 62153 58883
rect 58291 58502 60076 58697
rect 56099 58428 58005 58502
rect 53835 58424 55811 58428
rect 51760 58235 53551 58424
rect 47336 58125 51475 58235
rect 42800 58097 47025 58125
tri 42800 58010 42887 58097 ne
rect 42887 58010 47025 58097
tri 42600 57723 42887 58010 sw
tri 42887 57723 43174 58010 ne
rect 43174 57814 47025 58010
tri 47025 57814 47336 58125 sw
tri 47336 57814 47647 58125 ne
rect 47647 57950 51475 58125
tri 51475 57950 51760 58235 sw
tri 51760 57950 52045 58235 ne
rect 52045 58140 53551 58235
tri 53551 58140 53835 58424 sw
tri 53835 58140 54119 58424 ne
rect 54119 58140 55811 58424
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58332 58005 58428
tri 58005 58332 58175 58502 sw
tri 58291 58332 58461 58502 ne
rect 58461 58414 60076 58502
tri 60076 58414 60359 58697 sw
tri 60359 58414 60642 58697 ne
rect 60642 58600 62153 58697
tri 62153 58600 62436 58883 sw
tri 62436 58600 62719 58883 ne
rect 62719 58800 64212 58883
tri 64212 58800 64499 59087 sw
tri 64499 58800 64786 59087 ne
rect 64786 58920 70613 59087
rect 70669 58920 71000 60120
rect 64786 58800 71000 58920
rect 62719 58600 64499 58800
tri 64499 58600 64699 58800 sw
rect 60642 58414 62436 58600
rect 58461 58332 60359 58414
rect 56387 58140 58175 58332
rect 52045 57950 53835 58140
rect 47647 57814 51760 57950
rect 43174 57723 47336 57814
rect 41200 57436 42887 57723
tri 42887 57436 43174 57723 sw
tri 43174 57436 43461 57723 ne
rect 43461 57503 47336 57723
tri 47336 57503 47647 57814 sw
tri 47647 57503 47958 57814 ne
rect 47958 57665 51760 57814
tri 51760 57665 52045 57950 sw
tri 52045 57665 52330 57950 ne
rect 52330 57856 53835 57950
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 58048 56099 58140
tri 56099 58048 56191 58140 sw
tri 56387 58048 56479 58140 ne
rect 56479 58048 58175 58140
rect 54403 57856 56191 58048
rect 52330 57665 54119 57856
rect 47958 57503 52045 57665
rect 43461 57436 47647 57503
rect 41200 57430 43174 57436
tri 41200 57338 41292 57430 ne
rect 41292 57338 43174 57430
tri 41000 57138 41200 57338 sw
tri 41292 57138 41492 57338 ne
rect 41492 57321 43174 57338
tri 43174 57321 43289 57436 sw
tri 43461 57321 43576 57436 ne
rect 43576 57321 47647 57436
rect 41492 57138 43289 57321
rect 39600 56910 41200 57138
tri 41200 56910 41428 57138 sw
tri 41492 56910 41720 57138 ne
rect 41720 57034 43289 57138
tri 43289 57034 43576 57321 sw
tri 43576 57034 43863 57321 ne
rect 43863 57192 47647 57321
tri 47647 57192 47958 57503 sw
tri 47958 57192 48269 57503 ne
rect 48269 57395 52045 57503
tri 52045 57395 52315 57665 sw
tri 52330 57395 52600 57665 ne
rect 52600 57572 54119 57665
tri 54119 57572 54403 57856 sw
tri 54403 57572 54687 57856 ne
rect 54687 57760 56191 57856
tri 56191 57760 56479 58048 sw
tri 56479 57760 56767 58048 ne
rect 56767 58046 58175 58048
tri 58175 58046 58461 58332 sw
tri 58461 58046 58747 58332 ne
rect 58747 58131 60359 58332
tri 60359 58131 60642 58414 sw
tri 60642 58131 60925 58414 ne
rect 60925 58317 62436 58414
tri 62436 58317 62719 58600 sw
tri 62719 58317 63002 58600 ne
rect 63002 58317 71000 58600
rect 60925 58131 62719 58317
rect 58747 58046 60642 58131
rect 56767 57760 58461 58046
tri 58461 57760 58747 58046 sw
tri 58747 57760 59033 58046 ne
rect 59033 57946 60642 58046
tri 60642 57946 60827 58131 sw
tri 60925 57946 61110 58131 ne
rect 61110 58034 62719 58131
tri 62719 58034 63002 58317 sw
tri 63002 58034 63285 58317 ne
rect 63285 58034 71000 58317
rect 61110 57946 63002 58034
rect 59033 57760 60827 57946
rect 54687 57572 56479 57760
rect 52600 57395 54403 57572
rect 48269 57192 52315 57395
rect 43863 57034 47958 57192
rect 41720 56910 43576 57034
rect 39600 56758 41428 56910
tri 39600 56665 39693 56758 ne
rect 39693 56752 41428 56758
tri 41428 56752 41586 56910 sw
tri 41720 56752 41878 56910 ne
rect 41878 56752 43576 56910
rect 39693 56665 41586 56752
tri 39400 56465 39600 56665 sw
tri 39693 56465 39893 56665 ne
rect 39893 56465 41586 56665
rect 36400 56172 39600 56465
tri 39600 56172 39893 56465 sw
tri 39893 56172 40186 56465 ne
rect 40186 56460 41586 56465
tri 41586 56460 41878 56752 sw
tri 41878 56460 42170 56752 ne
rect 42170 56747 43576 56752
tri 43576 56747 43863 57034 sw
tri 43863 56747 44150 57034 ne
rect 44150 56910 47958 57034
tri 47958 56910 48240 57192 sw
tri 48269 56910 48551 57192 ne
rect 48551 57110 52315 57192
tri 52315 57110 52600 57395 sw
tri 52600 57110 52885 57395 ne
rect 52885 57288 54403 57395
tri 54403 57288 54687 57572 sw
tri 54687 57288 54971 57572 ne
rect 54971 57472 56479 57572
tri 56479 57472 56767 57760 sw
tri 56767 57472 57055 57760 ne
rect 57055 57666 58747 57760
tri 58747 57666 58841 57760 sw
tri 59033 57666 59127 57760 ne
rect 59127 57666 60827 57760
rect 57055 57472 58841 57666
rect 54971 57288 56767 57472
rect 52885 57110 54687 57288
rect 48551 56910 52600 57110
rect 44150 56803 48240 56910
tri 48240 56803 48347 56910 sw
tri 48551 56803 48658 56910 ne
rect 48658 56825 52600 56910
tri 52600 56825 52885 57110 sw
tri 52885 56825 53170 57110 ne
rect 53170 57108 54687 57110
tri 54687 57108 54867 57288 sw
tri 54971 57108 55151 57288 ne
rect 55151 57184 56767 57288
tri 56767 57184 57055 57472 sw
tri 57055 57184 57343 57472 ne
rect 57343 57380 58841 57472
tri 58841 57380 59127 57666 sw
tri 59127 57380 59413 57666 ne
rect 59413 57663 60827 57666
tri 60827 57663 61110 57946 sw
tri 61110 57663 61393 57946 ne
rect 61393 57766 63002 57946
tri 63002 57766 63270 58034 sw
tri 63285 57766 63553 58034 ne
rect 63553 57766 71000 58034
rect 61393 57663 63270 57766
rect 59413 57380 61110 57663
tri 61110 57380 61393 57663 sw
tri 61393 57380 61676 57663 ne
rect 61676 57483 63270 57663
tri 63270 57483 63553 57766 sw
tri 63553 57483 63836 57766 ne
rect 63836 57483 71000 57766
rect 61676 57380 63553 57483
rect 57343 57184 59127 57380
rect 55151 57108 57055 57184
rect 53170 56825 54867 57108
rect 48658 56803 52885 56825
rect 44150 56747 48347 56803
rect 42170 56460 43863 56747
tri 43863 56460 44150 56747 sw
tri 44150 56460 44437 56747 ne
rect 44437 56492 48347 56747
tri 48347 56492 48658 56803 sw
tri 48658 56492 48969 56803 ne
rect 48969 56540 52885 56803
tri 52885 56540 53170 56825 sw
tri 53170 56540 53455 56825 ne
rect 53455 56824 54867 56825
tri 54867 56824 55151 57108 sw
tri 55151 56824 55435 57108 ne
rect 55435 56896 57055 57108
tri 57055 56896 57343 57184 sw
tri 57343 56896 57631 57184 ne
rect 57631 57094 59127 57184
tri 59127 57094 59413 57380 sw
tri 59413 57094 59699 57380 ne
rect 59699 57283 61393 57380
tri 61393 57283 61490 57380 sw
tri 61676 57283 61773 57380 ne
rect 61773 57283 63553 57380
rect 59699 57094 61490 57283
rect 57631 56896 59413 57094
rect 55435 56824 57343 56896
rect 53455 56540 55151 56824
tri 55151 56540 55435 56824 sw
tri 55435 56540 55719 56824 ne
rect 55719 56736 57343 56824
tri 57343 56736 57503 56896 sw
tri 57631 56736 57791 56896 ne
rect 57791 56808 59413 56896
tri 59413 56808 59699 57094 sw
tri 59699 56808 59985 57094 ne
rect 59985 57000 61490 57094
tri 61490 57000 61773 57283 sw
tri 61773 57000 62056 57283 ne
rect 62056 57200 63553 57283
tri 63553 57200 63836 57483 sw
tri 63836 57200 64119 57483 ne
rect 64119 57200 71000 57483
rect 62056 57000 63836 57200
tri 63836 57000 64036 57200 sw
rect 59985 56808 61773 57000
rect 57791 56736 59699 56808
rect 55719 56540 57503 56736
rect 48969 56492 53170 56540
rect 44437 56460 48658 56492
rect 40186 56322 41878 56460
tri 41878 56322 42016 56460 sw
tri 42170 56322 42308 56460 ne
rect 42308 56322 44150 56460
rect 40186 56172 42016 56322
rect 36400 56145 39893 56172
tri 39893 56145 39920 56172 sw
tri 40186 56145 40213 56172 ne
rect 40213 56145 42016 56172
rect 36400 55852 39920 56145
tri 39920 55852 40213 56145 sw
tri 40213 55852 40506 56145 ne
rect 40506 56030 42016 56145
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56173 44150 56322
tri 44150 56173 44437 56460 sw
tri 44437 56173 44724 56460 ne
rect 44724 56181 48658 56460
tri 48658 56181 48969 56492 sw
tri 48969 56181 49280 56492 ne
rect 49280 56255 53170 56492
tri 53170 56255 53455 56540 sw
tri 53455 56255 53740 56540 ne
rect 53740 56444 55435 56540
tri 55435 56444 55531 56540 sw
tri 55719 56444 55815 56540 ne
rect 55815 56448 57503 56540
tri 57503 56448 57791 56736 sw
tri 57791 56448 58079 56736 ne
rect 58079 56522 59699 56736
tri 59699 56522 59985 56808 sw
tri 59985 56522 60271 56808 ne
rect 60271 56717 61773 56808
tri 61773 56717 62056 57000 sw
tri 62056 56717 62339 57000 ne
rect 62339 56910 71000 57000
rect 62339 56717 70613 56910
rect 60271 56522 62056 56717
rect 58079 56448 59985 56522
rect 55815 56444 57791 56448
rect 53740 56255 55531 56444
rect 49280 56181 53455 56255
rect 44724 56173 48969 56181
rect 42600 56030 44437 56173
rect 40506 55852 42308 56030
rect 36400 55559 40213 55852
tri 40213 55559 40506 55852 sw
tri 40506 55559 40799 55852 ne
rect 40799 55738 42308 55852
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55886 44437 56030
tri 44437 55886 44724 56173 sw
tri 44724 55886 45011 56173 ne
rect 45011 55886 48969 56173
rect 42892 55738 44724 55886
rect 40799 55559 42600 55738
rect 36400 55421 40506 55559
tri 36400 55324 36497 55421 ne
rect 36497 55324 40506 55421
tri 36200 55124 36400 55324 sw
tri 36497 55124 36697 55324 ne
rect 36697 55266 40506 55324
tri 40506 55266 40799 55559 sw
tri 40799 55266 41092 55559 ne
rect 41092 55446 42600 55559
tri 42600 55446 42892 55738 sw
tri 42892 55446 43184 55738 ne
rect 43184 55710 44724 55738
tri 44724 55710 44900 55886 sw
tri 45011 55710 45187 55886 ne
rect 45187 55870 48969 55886
tri 48969 55870 49280 56181 sw
tri 49280 55870 49591 56181 ne
rect 49591 55970 53455 56181
tri 53455 55970 53740 56255 sw
tri 53740 55970 54025 56255 ne
rect 54025 56160 55531 56255
tri 55531 56160 55815 56444 sw
tri 55815 56160 56099 56444 ne
rect 56099 56160 57791 56444
tri 57791 56160 58079 56448 sw
tri 58079 56160 58367 56448 ne
rect 58367 56352 59985 56448
tri 59985 56352 60155 56522 sw
tri 60271 56352 60441 56522 ne
rect 60441 56434 62056 56522
tri 62056 56434 62339 56717 sw
tri 62339 56434 62622 56717 ne
rect 62622 56434 70613 56717
rect 60441 56352 62339 56434
rect 58367 56160 60155 56352
rect 54025 55970 55815 56160
rect 49591 55870 53740 55970
rect 45187 55710 49280 55870
rect 43184 55559 44900 55710
tri 44900 55559 45051 55710 sw
tri 45187 55559 45338 55710 ne
rect 45338 55559 49280 55710
tri 49280 55559 49591 55870 sw
tri 49591 55559 49902 55870 ne
rect 49902 55685 53740 55870
tri 53740 55685 54025 55970 sw
tri 54025 55685 54310 55970 ne
rect 54310 55876 55815 55970
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 56068 58079 56160
tri 58079 56068 58171 56160 sw
tri 58367 56068 58459 56160 ne
rect 58459 56068 60155 56160
rect 56383 55876 58171 56068
rect 54310 55685 56099 55876
rect 49902 55559 54025 55685
rect 43184 55446 45051 55559
rect 41092 55266 42892 55446
rect 36697 55153 40799 55266
tri 40799 55153 40912 55266 sw
tri 41092 55153 41205 55266 ne
rect 41205 55154 42892 55266
tri 42892 55154 43184 55446 sw
tri 43184 55154 43476 55446 ne
rect 43476 55272 45051 55446
tri 45051 55272 45338 55559 sw
tri 45338 55272 45625 55559 ne
rect 45625 55272 49591 55559
rect 43476 55154 45338 55272
rect 41205 55153 43184 55154
rect 36697 55124 40912 55153
rect 33200 54827 36400 55124
tri 36400 54827 36697 55124 sw
tri 36697 54827 36994 55124 ne
rect 36994 54860 40912 55124
tri 40912 54860 41205 55153 sw
tri 41205 54860 41498 55153 ne
rect 41498 55064 43184 55153
tri 43184 55064 43274 55154 sw
tri 43476 55064 43566 55154 ne
rect 43566 55064 45338 55154
rect 41498 54860 43274 55064
rect 36994 54827 41205 54860
rect 33200 54674 36697 54827
tri 36697 54674 36850 54827 sw
tri 36994 54674 37147 54827 ne
rect 37147 54674 41205 54827
rect 33200 54377 36850 54674
tri 36850 54377 37147 54674 sw
tri 37147 54377 37444 54674 ne
rect 37444 54567 41205 54674
tri 41205 54567 41498 54860 sw
tri 41498 54567 41791 54860 ne
rect 41791 54772 43274 54860
tri 43274 54772 43566 55064 sw
tri 43566 54772 43858 55064 ne
rect 43858 55054 45338 55064
tri 45338 55054 45556 55272 sw
tri 45625 55054 45843 55272 ne
rect 45843 55248 49591 55272
tri 49591 55248 49902 55559 sw
tri 49902 55248 50213 55559 ne
rect 50213 55415 54025 55559
tri 54025 55415 54295 55685 sw
tri 54310 55415 54580 55685 ne
rect 54580 55592 56099 55685
tri 56099 55592 56383 55876 sw
tri 56383 55592 56667 55876 ne
rect 56667 55780 58171 55876
tri 58171 55780 58459 56068 sw
tri 58459 55780 58747 56068 ne
rect 58747 56066 60155 56068
tri 60155 56066 60441 56352 sw
tri 60441 56066 60727 56352 ne
rect 60727 56166 62339 56352
tri 62339 56166 62607 56434 sw
tri 62622 56166 62890 56434 ne
rect 62890 56166 70613 56434
rect 60727 56066 62607 56166
rect 58747 55780 60441 56066
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 55883 62607 56066
tri 62607 55883 62890 56166 sw
tri 62890 55883 63173 56166 ne
rect 63173 55883 70613 56166
rect 61013 55780 62890 55883
rect 56667 55592 58459 55780
rect 54580 55415 56383 55592
rect 50213 55248 54295 55415
rect 45843 55120 49902 55248
tri 49902 55120 50030 55248 sw
tri 50213 55120 50341 55248 ne
rect 50341 55130 54295 55248
tri 54295 55130 54580 55415 sw
tri 54580 55130 54865 55415 ne
rect 54865 55308 56383 55415
tri 56383 55308 56667 55592 sw
tri 56667 55308 56951 55592 ne
rect 56951 55492 58459 55592
tri 58459 55492 58747 55780 sw
tri 58747 55492 59035 55780 ne
rect 59035 55686 60727 55780
tri 60727 55686 60821 55780 sw
tri 61013 55686 61107 55780 ne
rect 61107 55686 62890 55780
rect 59035 55492 60821 55686
rect 56951 55308 58747 55492
rect 54865 55130 56667 55308
rect 50341 55120 54580 55130
rect 45843 55054 50030 55120
rect 43858 54772 45556 55054
rect 41791 54567 43566 54772
rect 37444 54377 41498 54567
rect 33200 54080 37147 54377
tri 37147 54080 37444 54377 sw
tri 37444 54080 37741 54377 ne
rect 37741 54274 41498 54377
tri 41498 54274 41791 54567 sw
tri 41791 54274 42084 54567 ne
rect 42084 54480 43566 54567
tri 43566 54480 43858 54772 sw
tri 43858 54480 44150 54772 ne
rect 44150 54767 45556 54772
tri 45556 54767 45843 55054 sw
tri 45843 54767 46130 55054 ne
rect 46130 54809 50030 55054
tri 50030 54809 50341 55120 sw
tri 50341 54809 50652 55120 ne
rect 50652 54845 54580 55120
tri 54580 54845 54865 55130 sw
tri 54865 54845 55150 55130 ne
rect 55150 55128 56667 55130
tri 56667 55128 56847 55308 sw
tri 56951 55128 57131 55308 ne
rect 57131 55204 58747 55308
tri 58747 55204 59035 55492 sw
tri 59035 55204 59323 55492 ne
rect 59323 55400 60821 55492
tri 60821 55400 61107 55686 sw
tri 61107 55400 61393 55686 ne
rect 61393 55600 62890 55686
tri 62890 55600 63173 55883 sw
tri 63173 55600 63456 55883 ne
rect 63456 55710 70613 55883
rect 70669 55710 71000 56910
rect 63456 55600 71000 55710
rect 61393 55400 63173 55600
tri 63173 55400 63373 55600 sw
rect 59323 55204 61107 55400
rect 57131 55128 59035 55204
rect 55150 54845 56847 55128
rect 50652 54809 54865 54845
rect 46130 54767 50341 54809
rect 44150 54480 45843 54767
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54498 50341 54767
tri 50341 54498 50652 54809 sw
tri 50652 54498 50963 54809 ne
rect 50963 54560 54865 54809
tri 54865 54560 55150 54845 sw
tri 55150 54560 55435 54845 ne
rect 55435 54844 56847 54845
tri 56847 54844 57131 55128 sw
tri 57131 54844 57415 55128 ne
rect 57415 54916 59035 55128
tri 59035 54916 59323 55204 sw
tri 59323 54916 59611 55204 ne
rect 59611 55114 61107 55204
tri 61107 55114 61393 55400 sw
tri 61393 55114 61679 55400 ne
rect 61679 55302 71000 55400
rect 61679 55114 70613 55302
rect 59611 54916 61393 55114
rect 57415 54844 59323 54916
rect 55435 54560 57131 54844
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54756 59323 54844
tri 59323 54756 59483 54916 sw
tri 59611 54756 59771 54916 ne
rect 59771 54828 61393 54916
tri 61393 54828 61679 55114 sw
tri 61679 54828 61965 55114 ne
rect 61965 54828 70613 55114
rect 59771 54756 61679 54828
rect 57699 54560 59483 54756
rect 50963 54498 55150 54560
rect 46417 54480 50652 54498
rect 42084 54274 43858 54480
rect 37741 54080 41791 54274
tri 33200 53992 33288 54080 ne
rect 33288 53992 37444 54080
tri 33000 53792 33200 53992 sw
tri 33288 53792 33488 53992 ne
rect 33488 53792 37444 53992
rect 30000 53504 33200 53792
tri 33200 53504 33488 53792 sw
tri 33488 53504 33776 53792 ne
rect 33776 53783 37444 53792
tri 37444 53783 37741 54080 sw
tri 37741 53783 38038 54080 ne
rect 38038 53981 41791 54080
tri 41791 53981 42084 54274 sw
tri 42084 53981 42377 54274 ne
rect 42377 54188 43858 54274
tri 43858 54188 44150 54480 sw
tri 44150 54188 44442 54480 ne
rect 44442 54193 46130 54480
tri 46130 54193 46417 54480 sw
tri 46417 54193 46704 54480 ne
rect 46704 54193 50652 54480
rect 44442 54188 46417 54193
rect 42377 53981 44150 54188
rect 38038 53783 42084 53981
rect 33776 53673 37741 53783
tri 37741 53673 37851 53783 sw
tri 38038 53673 38148 53783 ne
rect 38148 53722 42084 53783
tri 42084 53722 42343 53981 sw
tri 42377 53722 42636 53981 ne
rect 42636 53896 44150 53981
tri 44150 53896 44442 54188 sw
tri 44442 53896 44734 54188 ne
rect 44734 53906 46417 54188
tri 46417 53906 46704 54193 sw
tri 46704 53906 46991 54193 ne
rect 46991 54187 50652 54193
tri 50652 54187 50963 54498 sw
tri 50963 54187 51274 54498 ne
rect 51274 54275 55150 54498
tri 55150 54275 55435 54560 sw
tri 55435 54275 55720 54560 ne
rect 55720 54464 57415 54560
tri 57415 54464 57511 54560 sw
tri 57699 54464 57795 54560 ne
rect 57795 54468 59483 54560
tri 59483 54468 59771 54756 sw
tri 59771 54468 60059 54756 ne
rect 60059 54572 61679 54756
tri 61679 54572 61935 54828 sw
tri 61965 54572 62221 54828 ne
rect 62221 54572 70613 54828
rect 60059 54468 61935 54572
rect 57795 54464 59771 54468
rect 55720 54275 57511 54464
rect 51274 54187 55435 54275
rect 46991 53906 50963 54187
rect 44734 53896 46704 53906
rect 42636 53722 44442 53896
rect 38148 53673 42343 53722
rect 33776 53504 37851 53673
rect 30000 53216 33488 53504
tri 33488 53216 33776 53504 sw
tri 33776 53216 34064 53504 ne
rect 34064 53376 37851 53504
tri 37851 53376 38148 53673 sw
tri 38148 53376 38445 53673 ne
rect 38445 53466 42343 53673
tri 42343 53466 42599 53722 sw
tri 42636 53466 42892 53722 ne
rect 42892 53604 44442 53722
tri 44442 53604 44734 53896 sw
tri 44734 53604 45026 53896 ne
rect 45026 53619 46704 53896
tri 46704 53619 46991 53906 sw
tri 46991 53619 47278 53906 ne
rect 47278 53876 50963 53906
tri 50963 53876 51274 54187 sw
tri 51274 53876 51585 54187 ne
rect 51585 53990 55435 54187
tri 55435 53990 55720 54275 sw
tri 55720 53990 56005 54275 ne
rect 56005 54180 57511 54275
tri 57511 54180 57795 54464 sw
tri 57795 54180 58079 54464 ne
rect 58079 54180 59771 54464
tri 59771 54180 60059 54468 sw
tri 60059 54180 60347 54468 ne
rect 60347 54286 61935 54468
tri 61935 54286 62221 54572 sw
tri 62221 54286 62507 54572 ne
rect 62507 54286 70613 54572
rect 60347 54180 62221 54286
rect 56005 53990 57795 54180
rect 51585 53876 55720 53990
rect 47278 53619 51274 53876
rect 45026 53604 46991 53619
rect 42892 53466 44734 53604
rect 38445 53376 42599 53466
rect 34064 53216 38148 53376
rect 30000 52928 33776 53216
tri 33776 52928 34064 53216 sw
tri 34064 52928 34352 53216 ne
rect 34352 53079 38148 53216
tri 38148 53079 38445 53376 sw
tri 38445 53079 38742 53376 ne
rect 38742 53173 42599 53376
tri 42599 53173 42892 53466 sw
tri 42892 53173 43185 53466 ne
rect 43185 53464 44734 53466
tri 44734 53464 44874 53604 sw
tri 45026 53464 45166 53604 ne
rect 45166 53464 46991 53604
rect 43185 53173 44874 53464
rect 38742 53079 42892 53173
rect 34352 52928 38445 53079
rect 30000 52748 34064 52928
tri 30000 52654 30094 52748 ne
rect 30094 52654 34064 52748
tri 29800 52454 30000 52654 sw
tri 30094 52454 30294 52654 ne
rect 30294 52640 34064 52654
tri 34064 52640 34352 52928 sw
tri 34352 52640 34640 52928 ne
rect 34640 52782 38445 52928
tri 38445 52782 38742 53079 sw
tri 38742 52782 39039 53079 ne
rect 39039 52880 42892 53079
tri 42892 52880 43185 53173 sw
tri 43185 52880 43478 53173 ne
rect 43478 53172 44874 53173
tri 44874 53172 45166 53464 sw
tri 45166 53172 45458 53464 ne
rect 45458 53361 46991 53464
tri 46991 53361 47249 53619 sw
tri 47278 53361 47536 53619 ne
rect 47536 53565 51274 53619
tri 51274 53565 51585 53876 sw
tri 51585 53565 51896 53876 ne
rect 51896 53705 55720 53876
tri 55720 53705 56005 53990 sw
tri 56005 53705 56290 53990 ne
rect 56290 53896 57795 53990
tri 57795 53896 58079 54180 sw
tri 58079 53896 58363 54180 ne
rect 58363 54088 60059 54180
tri 60059 54088 60151 54180 sw
tri 60347 54088 60439 54180 ne
rect 60439 54088 62221 54180
rect 58363 53896 60151 54088
rect 56290 53705 58079 53896
rect 51896 53565 56005 53705
rect 47536 53361 51585 53565
rect 45458 53172 47249 53361
rect 43478 52880 45166 53172
tri 45166 52880 45458 53172 sw
tri 45458 52880 45750 53172 ne
rect 45750 53074 47249 53172
tri 47249 53074 47536 53361 sw
tri 47536 53074 47823 53361 ne
rect 47823 53254 51585 53361
tri 51585 53254 51896 53565 sw
tri 51896 53254 52207 53565 ne
rect 52207 53435 56005 53565
tri 56005 53435 56275 53705 sw
tri 56290 53435 56560 53705 ne
rect 56560 53612 58079 53705
tri 58079 53612 58363 53896 sw
tri 58363 53612 58647 53896 ne
rect 58647 53800 60151 53896
tri 60151 53800 60439 54088 sw
tri 60439 53800 60727 54088 ne
rect 60727 54000 62221 54088
tri 62221 54000 62507 54286 sw
tri 62507 54000 62793 54286 ne
rect 62793 54102 70613 54286
rect 70669 54102 71000 55302
rect 62793 54000 71000 54102
rect 60727 53800 62507 54000
tri 62507 53800 62707 54000 sw
rect 58647 53612 60439 53800
rect 56560 53435 58363 53612
rect 52207 53254 56275 53435
rect 47823 53074 51896 53254
rect 45750 52880 47536 53074
rect 39039 52782 43185 52880
rect 34640 52640 38742 52782
rect 30294 52454 34352 52640
rect 26800 52160 30000 52454
tri 30000 52160 30294 52454 sw
tri 30294 52160 30588 52454 ne
rect 30588 52372 34352 52454
tri 34352 52372 34620 52640 sw
tri 34640 52372 34908 52640 ne
rect 34908 52485 38742 52640
tri 38742 52485 39039 52782 sw
tri 39039 52485 39336 52782 ne
rect 39336 52587 43185 52782
tri 43185 52587 43478 52880 sw
tri 43478 52587 43771 52880 ne
rect 43771 52804 45458 52880
tri 45458 52804 45534 52880 sw
tri 45750 52804 45826 52880 ne
rect 45826 52804 47536 52880
rect 43771 52587 45534 52804
rect 39336 52485 43478 52587
rect 34908 52372 39039 52485
rect 30588 52160 34620 52372
rect 26800 51998 30294 52160
tri 30294 51998 30456 52160 sw
tri 30588 51998 30750 52160 ne
rect 30750 52084 34620 52160
tri 34620 52084 34908 52372 sw
tri 34908 52084 35196 52372 ne
rect 35196 52188 39039 52372
tri 39039 52188 39336 52485 sw
tri 39336 52188 39633 52485 ne
rect 39633 52294 43478 52485
tri 43478 52294 43771 52587 sw
tri 43771 52294 44064 52587 ne
rect 44064 52512 45534 52587
tri 45534 52512 45826 52804 sw
tri 45826 52512 46118 52804 ne
rect 46118 52787 47536 52804
tri 47536 52787 47823 53074 sw
tri 47823 52787 48110 53074 ne
rect 48110 52943 51896 53074
tri 51896 52943 52207 53254 sw
tri 52207 52943 52518 53254 ne
rect 52518 53150 56275 53254
tri 56275 53150 56560 53435 sw
tri 56560 53150 56845 53435 ne
rect 56845 53328 58363 53435
tri 58363 53328 58647 53612 sw
tri 58647 53328 58931 53612 ne
rect 58931 53512 60439 53612
tri 60439 53512 60727 53800 sw
tri 60727 53512 61015 53800 ne
rect 61015 53722 71000 53800
rect 61015 53512 70613 53722
rect 58931 53328 60727 53512
rect 56845 53150 58647 53328
rect 52518 52943 56560 53150
rect 48110 52861 52207 52943
tri 52207 52861 52289 52943 sw
tri 52518 52861 52600 52943 ne
rect 52600 52865 56560 52943
tri 56560 52865 56845 53150 sw
tri 56845 52865 57130 53150 ne
rect 57130 53148 58647 53150
tri 58647 53148 58827 53328 sw
tri 58931 53148 59111 53328 ne
rect 59111 53224 60727 53328
tri 60727 53224 61015 53512 sw
tri 61015 53224 61303 53512 ne
rect 61303 53224 70613 53512
rect 59111 53148 61015 53224
rect 57130 52865 58827 53148
rect 52600 52861 56845 52865
rect 48110 52787 52289 52861
rect 46118 52512 47823 52787
rect 44064 52500 45826 52512
tri 45826 52500 45838 52512 sw
tri 46118 52500 46130 52512 ne
rect 46130 52500 47823 52512
tri 47823 52500 48110 52787 sw
tri 48110 52500 48397 52787 ne
rect 48397 52550 52289 52787
tri 52289 52550 52600 52861 sw
tri 52600 52550 52911 52861 ne
rect 52911 52580 56845 52861
tri 56845 52580 57130 52865 sw
tri 57130 52580 57415 52865 ne
rect 57415 52864 58827 52865
tri 58827 52864 59111 53148 sw
tri 59111 52864 59395 53148 ne
rect 59395 52976 61015 53148
tri 61015 52976 61263 53224 sw
tri 61303 52976 61551 53224 ne
rect 61551 52976 70613 53224
rect 59395 52864 61263 52976
rect 57415 52580 59111 52864
tri 59111 52580 59395 52864 sw
tri 59395 52580 59679 52864 ne
rect 59679 52688 61263 52864
tri 61263 52688 61551 52976 sw
tri 61551 52688 61839 52976 ne
rect 61839 52688 70613 52976
rect 59679 52580 61551 52688
rect 52911 52550 57130 52580
rect 48397 52500 52600 52550
rect 44064 52294 45838 52500
rect 39633 52188 43771 52294
rect 35196 52084 39336 52188
rect 30750 51998 34908 52084
rect 26800 51704 30456 51998
tri 30456 51704 30750 51998 sw
tri 30750 51704 31044 51998 ne
rect 31044 51796 34908 51998
tri 34908 51796 35196 52084 sw
tri 35196 51796 35484 52084 ne
rect 35484 51891 39336 52084
tri 39336 51891 39633 52188 sw
tri 39633 51891 39930 52188 ne
rect 39930 52001 43771 52188
tri 43771 52001 44064 52294 sw
tri 44064 52001 44357 52294 ne
rect 44357 52208 45838 52294
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52213 48110 52500
tri 48110 52213 48397 52500 sw
tri 48397 52213 48684 52500 ne
rect 48684 52239 52600 52500
tri 52600 52239 52911 52550 sw
tri 52911 52239 53222 52550 ne
rect 53222 52295 57130 52550
tri 57130 52295 57415 52580 sw
tri 57415 52295 57700 52580 ne
rect 57700 52484 59395 52580
tri 59395 52484 59491 52580 sw
tri 59679 52484 59775 52580 ne
rect 59775 52484 61551 52580
rect 57700 52295 59491 52484
rect 53222 52239 57415 52295
rect 48684 52213 52911 52239
rect 46422 52208 48397 52213
rect 44357 52001 46130 52208
rect 39930 51891 44064 52001
rect 35484 51796 39633 51891
rect 31044 51704 35196 51796
rect 26800 51410 30750 51704
tri 30750 51410 31044 51704 sw
tri 31044 51410 31338 51704 ne
rect 31338 51508 35196 51704
tri 35196 51508 35484 51796 sw
tri 35484 51508 35772 51796 ne
rect 35772 51661 39633 51796
tri 39633 51661 39863 51891 sw
tri 39930 51661 40160 51891 ne
rect 40160 51779 44064 51891
tri 44064 51779 44286 52001 sw
tri 44357 51779 44579 52001 ne
rect 44579 51916 46130 52001
tri 46130 51916 46422 52208 sw
tri 46422 51916 46714 52208 ne
rect 46714 51926 48397 52208
tri 48397 51926 48684 52213 sw
tri 48684 51926 48971 52213 ne
rect 48971 51928 52911 52213
tri 52911 51928 53222 52239 sw
tri 53222 51928 53533 52239 ne
rect 53533 52010 57415 52239
tri 57415 52010 57700 52295 sw
tri 57700 52010 57985 52295 ne
rect 57985 52200 59491 52295
tri 59491 52200 59775 52484 sw
tri 59775 52200 60059 52484 ne
rect 60059 52400 61551 52484
tri 61551 52400 61839 52688 sw
tri 61839 52400 62127 52688 ne
rect 62127 52522 70613 52688
rect 70669 52522 71000 53722
rect 62127 52400 71000 52522
rect 60059 52200 61839 52400
tri 61839 52200 62039 52400 sw
rect 57985 52010 59775 52200
rect 53533 51928 57700 52010
rect 48971 51926 53222 51928
rect 46714 51916 48684 51926
rect 44579 51779 46422 51916
rect 40160 51661 44286 51779
rect 35772 51508 39863 51661
rect 31338 51410 35484 51508
tri 26800 51320 26890 51410 ne
rect 26890 51320 31044 51410
tri 26600 51220 26700 51320 sw
tri 26890 51220 26990 51320 ne
rect 26990 51220 31044 51320
tri 31044 51220 31234 51410 sw
tri 31338 51220 31528 51410 ne
rect 31528 51220 35484 51410
tri 35484 51220 35772 51508 sw
tri 35772 51220 36060 51508 ne
rect 36060 51364 39863 51508
tri 39863 51364 40160 51661 sw
tri 40160 51364 40457 51661 ne
rect 40457 51486 44286 51661
tri 44286 51486 44579 51779 sw
tri 44579 51486 44872 51779 ne
rect 44872 51624 46422 51779
tri 46422 51624 46714 51916 sw
tri 46714 51624 47006 51916 ne
rect 47006 51880 48684 51916
tri 48684 51880 48730 51926 sw
tri 48971 51880 49017 51926 ne
rect 49017 51880 53222 51926
rect 47006 51624 48730 51880
rect 44872 51486 46714 51624
rect 40457 51364 44579 51486
rect 36060 51220 40160 51364
rect 25200 50930 26700 51220
tri 26700 50930 26990 51220 sw
tri 26990 50930 27280 51220 ne
rect 27280 50930 31234 51220
rect 25200 50740 26990 50930
tri 25200 50651 25289 50740 ne
rect 25289 50651 26990 50740
tri 25000 50451 25200 50651 sw
tri 25289 50451 25489 50651 ne
rect 25489 50650 26990 50651
tri 26990 50650 27270 50930 sw
tri 27280 50650 27560 50930 ne
rect 27560 50926 31234 50930
tri 31234 50926 31528 51220 sw
tri 31528 50926 31822 51220 ne
rect 31822 50932 35772 51220
tri 35772 50932 36060 51220 sw
tri 36060 50932 36348 51220 ne
rect 36348 51067 40160 51220
tri 40160 51067 40457 51364 sw
tri 40457 51067 40754 51364 ne
rect 40754 51193 44579 51364
tri 44579 51193 44872 51486 sw
tri 44872 51193 45165 51486 ne
rect 45165 51484 46714 51486
tri 46714 51484 46854 51624 sw
tri 47006 51484 47146 51624 ne
rect 47146 51593 48730 51624
tri 48730 51593 49017 51880 sw
tri 49017 51593 49304 51880 ne
rect 49304 51617 53222 51880
tri 53222 51617 53533 51928 sw
tri 53533 51617 53844 51928 ne
rect 53844 51725 57700 51928
tri 57700 51725 57985 52010 sw
tri 57985 51725 58270 52010 ne
rect 58270 51916 59775 52010
tri 59775 51916 60059 52200 sw
tri 60059 51916 60343 52200 ne
rect 60343 51916 71000 52200
rect 58270 51725 60059 51916
rect 53844 51617 57985 51725
rect 49304 51593 53533 51617
rect 47146 51484 49017 51593
rect 45165 51193 46854 51484
rect 40754 51067 44872 51193
rect 36348 50932 40457 51067
rect 31822 50926 36060 50932
rect 27560 50650 31528 50926
rect 25489 50451 27270 50650
rect 23600 50360 25200 50451
tri 25200 50360 25291 50451 sw
tri 25489 50360 25580 50451 ne
rect 25580 50360 27270 50451
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50632 31528 50650
tri 31528 50632 31822 50926 sw
tri 31822 50632 32116 50926 ne
rect 32116 50752 36060 50926
tri 36060 50752 36240 50932 sw
tri 36348 50752 36528 50932 ne
rect 36528 50770 40457 50932
tri 40457 50770 40754 51067 sw
tri 40754 50770 41051 51067 ne
rect 41051 50900 44872 51067
tri 44872 50900 45165 51193 sw
tri 45165 50900 45458 51193 ne
rect 45458 51192 46854 51193
tri 46854 51192 47146 51484 sw
tri 47146 51192 47438 51484 ne
rect 47438 51306 49017 51484
tri 49017 51306 49304 51593 sw
tri 49304 51306 49591 51593 ne
rect 49591 51306 53533 51593
tri 53533 51306 53844 51617 sw
tri 53844 51306 54155 51617 ne
rect 54155 51455 57985 51617
tri 57985 51455 58255 51725 sw
tri 58270 51455 58540 51725 ne
rect 58540 51632 60059 51725
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58540 51455 60343 51632
rect 54155 51306 58255 51455
rect 47438 51192 49304 51306
rect 45458 50900 47146 51192
tri 47146 50900 47438 51192 sw
tri 47438 50900 47730 51192 ne
rect 47730 51019 49304 51192
tri 49304 51019 49591 51306 sw
tri 49591 51019 49878 51306 ne
rect 49878 51019 53844 51306
rect 47730 50900 49591 51019
rect 41051 50770 45165 50900
rect 36528 50752 40754 50770
rect 32116 50632 36240 50752
rect 27850 50360 31822 50632
rect 23600 50071 25291 50360
tri 25291 50071 25580 50360 sw
tri 25580 50071 25869 50360 ne
rect 25869 50071 27560 50360
tri 23600 49974 23697 50071 ne
rect 23697 49974 25580 50071
tri 23400 49774 23600 49974 sw
tri 23697 49774 23897 49974 ne
rect 23897 49918 25580 49974
tri 25580 49918 25733 50071 sw
tri 25869 49918 26022 50071 ne
rect 26022 50070 27560 50071
tri 27560 50070 27850 50360 sw
tri 27850 50070 28140 50360 ne
rect 28140 50338 31822 50360
tri 31822 50338 32116 50632 sw
tri 32116 50338 32410 50632 ne
rect 32410 50464 36240 50632
tri 36240 50464 36528 50752 sw
tri 36528 50464 36816 50752 ne
rect 36816 50473 40754 50752
tri 40754 50473 41051 50770 sw
tri 41051 50473 41348 50770 ne
rect 41348 50607 45165 50770
tri 45165 50607 45458 50900 sw
tri 45458 50607 45751 50900 ne
rect 45751 50812 47438 50900
tri 47438 50812 47526 50900 sw
tri 47730 50812 47818 50900 ne
rect 47818 50812 49591 50900
rect 45751 50607 47526 50812
rect 41348 50473 45458 50607
rect 36816 50464 41051 50473
rect 32410 50338 36528 50464
rect 28140 50070 32116 50338
rect 26022 49974 27850 50070
tri 27850 49974 27946 50070 sw
tri 28140 49974 28236 50070 ne
rect 28236 50044 32116 50070
tri 32116 50044 32410 50338 sw
tri 32410 50044 32704 50338 ne
rect 32704 50176 36528 50338
tri 36528 50176 36816 50464 sw
tri 36816 50176 37104 50464 ne
rect 37104 50176 41051 50464
tri 41051 50176 41348 50473 sw
tri 41348 50176 41645 50473 ne
rect 41645 50314 45458 50473
tri 45458 50314 45751 50607 sw
tri 45751 50314 46044 50607 ne
rect 46044 50520 47526 50607
tri 47526 50520 47818 50812 sw
tri 47818 50520 48110 50812 ne
rect 48110 50807 49591 50812
tri 49591 50807 49803 51019 sw
tri 49878 50807 50090 51019 ne
rect 50090 50995 53844 51019
tri 53844 50995 54155 51306 sw
tri 54155 50995 54466 51306 ne
rect 54466 51170 58255 51306
tri 58255 51170 58540 51455 sw
tri 58540 51170 58825 51455 ne
rect 58825 51368 60343 51455
tri 60343 51368 60607 51632 sw
tri 60627 51368 60891 51632 ne
rect 60891 51368 71000 51632
rect 58825 51170 60607 51368
rect 54466 50995 58540 51170
rect 50090 50871 54155 50995
tri 54155 50871 54279 50995 sw
tri 54466 50871 54590 50995 ne
rect 54590 50885 58540 50995
tri 58540 50885 58825 51170 sw
tri 58825 50885 59110 51170 ne
rect 59110 51084 60607 51170
tri 60607 51084 60891 51368 sw
tri 60891 51084 61175 51368 ne
rect 61175 51084 71000 51368
rect 59110 50885 60891 51084
rect 54590 50871 58825 50885
rect 50090 50807 54279 50871
rect 48110 50520 49803 50807
tri 49803 50520 50090 50807 sw
tri 50090 50520 50377 50807 ne
rect 50377 50560 54279 50807
tri 54279 50560 54590 50871 sw
tri 54590 50560 54901 50871 ne
rect 54901 50600 58825 50871
tri 58825 50600 59110 50885 sw
tri 59110 50600 59395 50885 ne
rect 59395 50800 60891 50885
tri 60891 50800 61175 51084 sw
tri 61175 50800 61459 51084 ne
rect 61459 50800 71000 51084
rect 59395 50600 61175 50800
tri 61175 50600 61375 50800 sw
rect 54901 50560 59110 50600
rect 50377 50520 54590 50560
rect 46044 50314 47818 50520
rect 41645 50176 45751 50314
rect 32704 50044 36816 50176
rect 28236 49974 32410 50044
rect 26022 49918 27946 49974
rect 23897 49774 25733 49918
rect 20400 49477 23600 49774
tri 23600 49477 23897 49774 sw
tri 23897 49477 24194 49774 ne
rect 24194 49629 25733 49774
tri 25733 49629 26022 49918 sw
tri 26022 49629 26311 49918 ne
rect 26311 49684 27946 49918
tri 27946 49684 28236 49974 sw
tri 28236 49684 28526 49974 ne
rect 28526 49750 32410 49974
tri 32410 49750 32704 50044 sw
tri 32704 49750 32998 50044 ne
rect 32998 49888 36816 50044
tri 36816 49888 37104 50176 sw
tri 37104 49888 37392 50176 ne
rect 37392 49888 41348 50176
rect 32998 49750 37104 49888
rect 28526 49684 32704 49750
rect 26311 49629 28236 49684
rect 24194 49477 26022 49629
rect 20400 49354 23897 49477
tri 23897 49354 24020 49477 sw
tri 24194 49354 24317 49477 ne
rect 24317 49354 26022 49477
rect 20400 49057 24020 49354
tri 24020 49057 24317 49354 sw
tri 24317 49057 24614 49354 ne
rect 24614 49340 26022 49354
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49394 28236 49629
tri 28236 49394 28526 49684 sw
tri 28526 49394 28816 49684 ne
rect 28816 49490 32704 49684
tri 32704 49490 32964 49750 sw
tri 32998 49490 33258 49750 ne
rect 33258 49600 37104 49750
tri 37104 49600 37392 49888 sw
tri 37392 49600 37680 49888 ne
rect 37680 49879 41348 49888
tri 41348 49879 41645 50176 sw
tri 41645 49879 41942 50176 ne
rect 41942 50021 45751 50176
tri 45751 50021 46044 50314 sw
tri 46044 50021 46337 50314 ne
rect 46337 50228 47818 50314
tri 47818 50228 48110 50520 sw
tri 48110 50228 48402 50520 ne
rect 48402 50249 50090 50520
tri 50090 50249 50361 50520 sw
tri 50377 50249 50648 50520 ne
rect 50648 50249 54590 50520
tri 54590 50249 54901 50560 sw
tri 54901 50249 55212 50560 ne
rect 55212 50315 59110 50560
tri 59110 50315 59395 50600 sw
tri 59395 50315 59680 50600 ne
rect 59680 50315 71000 50600
rect 55212 50249 59395 50315
rect 48402 50228 50361 50249
rect 46337 50021 48110 50228
rect 41942 49879 46044 50021
rect 37680 49726 41645 49879
tri 41645 49726 41798 49879 sw
tri 41942 49726 42095 49879 ne
rect 42095 49799 46044 49879
tri 46044 49799 46266 50021 sw
tri 46337 49799 46559 50021 ne
rect 46559 49936 48110 50021
tri 48110 49936 48402 50228 sw
tri 48402 49936 48694 50228 ne
rect 48694 49962 50361 50228
tri 50361 49962 50648 50249 sw
tri 50648 49962 50935 50249 ne
rect 50935 49962 54901 50249
rect 48694 49936 50648 49962
rect 46559 49799 48402 49936
rect 42095 49726 46266 49799
rect 37680 49600 41798 49726
rect 33258 49490 37392 49600
rect 28816 49394 32964 49490
rect 26600 49340 28526 49394
rect 24614 49057 26311 49340
rect 20400 48760 24317 49057
tri 24317 48760 24614 49057 sw
tri 24614 48760 24911 49057 ne
rect 24911 49051 26311 49057
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49250 28526 49340
tri 28526 49250 28670 49394 sw
tri 28816 49250 28960 49394 ne
rect 28960 49250 32964 49394
rect 26889 49051 28670 49250
rect 24911 48762 26600 49051
tri 26600 48762 26889 49051 sw
tri 26889 48762 27178 49051 ne
rect 27178 48960 28670 49051
tri 28670 48960 28960 49250 sw
tri 28960 48960 29250 49250 ne
rect 29250 49196 32964 49250
tri 32964 49196 33258 49490 sw
tri 33258 49196 33552 49490 ne
rect 33552 49312 37392 49490
tri 37392 49312 37680 49600 sw
tri 37680 49312 37968 49600 ne
rect 37968 49429 41798 49600
tri 41798 49429 42095 49726 sw
tri 42095 49429 42392 49726 ne
rect 42392 49506 46266 49726
tri 46266 49506 46559 49799 sw
tri 46559 49506 46852 49799 ne
rect 46852 49644 48402 49799
tri 48402 49644 48694 49936 sw
tri 48694 49644 48986 49936 ne
rect 48986 49675 50648 49936
tri 50648 49675 50935 49962 sw
tri 50935 49675 51222 49962 ne
rect 51222 49938 54901 49962
tri 54901 49938 55212 50249 sw
tri 55212 49938 55523 50249 ne
rect 55523 50030 59395 50249
tri 59395 50030 59680 50315 sw
tri 59680 50030 59965 50315 ne
rect 59965 50030 71000 50315
rect 55523 49938 59680 50030
rect 51222 49675 55212 49938
rect 48986 49644 50935 49675
rect 46852 49506 48694 49644
rect 42392 49429 46559 49506
rect 37968 49312 42095 49429
rect 33552 49196 37680 49312
rect 29250 48960 33258 49196
rect 27178 48762 28960 48960
rect 24911 48760 26889 48762
rect 20400 48730 24614 48760
tri 20400 48648 20482 48730 ne
rect 20482 48671 24614 48730
tri 24614 48671 24703 48760 sw
tri 24911 48671 25000 48760 ne
rect 25000 48671 26889 48760
rect 20482 48648 24703 48671
tri 20200 48448 20400 48648 sw
tri 20482 48448 20682 48648 ne
rect 20682 48448 24703 48648
rect 17200 48166 20400 48448
tri 20400 48166 20682 48448 sw
tri 20682 48166 20964 48448 ne
rect 20964 48374 24703 48448
tri 24703 48374 25000 48671 sw
tri 25000 48374 25297 48671 ne
rect 25297 48669 26889 48671
tri 26889 48669 26982 48762 sw
tri 27178 48669 27271 48762 ne
rect 27271 48670 28960 48762
tri 28960 48670 29250 48960 sw
tri 29250 48670 29540 48960 ne
rect 29540 48902 33258 48960
tri 33258 48902 33552 49196 sw
tri 33552 48902 33846 49196 ne
rect 33846 49024 37680 49196
tri 37680 49024 37968 49312 sw
tri 37968 49024 38256 49312 ne
rect 38256 49132 42095 49312
tri 42095 49132 42392 49429 sw
tri 42392 49132 42689 49429 ne
rect 42689 49213 46559 49429
tri 46559 49213 46852 49506 sw
tri 46852 49213 47145 49506 ne
rect 47145 49504 48694 49506
tri 48694 49504 48834 49644 sw
tri 48986 49504 49126 49644 ne
rect 49126 49504 50935 49644
rect 47145 49213 48834 49504
rect 42689 49132 46852 49213
rect 38256 49024 42392 49132
rect 33846 48902 37968 49024
rect 29540 48670 33552 48902
rect 27271 48669 29250 48670
rect 25297 48380 26982 48669
tri 26982 48380 27271 48669 sw
tri 27271 48380 27560 48669 ne
rect 27560 48380 29250 48669
tri 29250 48380 29540 48670 sw
tri 29540 48380 29830 48670 ne
rect 29830 48608 33552 48670
tri 33552 48608 33846 48902 sw
tri 33846 48608 34140 48902 ne
rect 34140 48736 37968 48902
tri 37968 48736 38256 49024 sw
tri 38256 48736 38544 49024 ne
rect 38544 48835 42392 49024
tri 42392 48835 42689 49132 sw
tri 42689 48835 42986 49132 ne
rect 42986 48920 46852 49132
tri 46852 48920 47145 49213 sw
tri 47145 48920 47438 49213 ne
rect 47438 49212 48834 49213
tri 48834 49212 49126 49504 sw
tri 49126 49212 49418 49504 ne
rect 49418 49419 50935 49504
tri 50935 49419 51191 49675 sw
tri 51222 49419 51478 49675 ne
rect 51478 49627 55212 49675
tri 55212 49627 55523 49938 sw
tri 55523 49627 55834 49938 ne
rect 55834 49770 59680 49938
tri 59680 49770 59940 50030 sw
tri 59965 49770 60225 50030 ne
rect 60225 49770 71000 50030
rect 55834 49627 59940 49770
rect 51478 49419 55523 49627
rect 49418 49212 51191 49419
rect 47438 48920 49126 49212
tri 49126 48920 49418 49212 sw
tri 49418 48920 49710 49212 ne
rect 49710 49132 51191 49212
tri 51191 49132 51478 49419 sw
tri 51478 49132 51765 49419 ne
rect 51765 49316 55523 49419
tri 55523 49316 55834 49627 sw
tri 55834 49316 56145 49627 ne
rect 56145 49485 59940 49627
tri 59940 49485 60225 49770 sw
tri 60225 49485 60510 49770 ne
rect 60510 49485 71000 49770
rect 56145 49316 60225 49485
rect 51765 49132 55834 49316
rect 49710 48920 51478 49132
rect 42986 48835 47145 48920
rect 38544 48736 42689 48835
rect 34140 48608 38256 48736
rect 29830 48380 33846 48608
rect 25297 48374 27271 48380
rect 20964 48166 25000 48374
rect 17200 47884 20682 48166
tri 20682 47884 20964 48166 sw
tri 20964 47884 21246 48166 ne
rect 21246 48077 25000 48166
tri 25000 48077 25297 48374 sw
tri 25297 48077 25594 48374 ne
rect 25594 48091 27271 48374
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48091 29540 48380
rect 25594 48077 27560 48091
rect 21246 47884 25297 48077
rect 17200 47602 20964 47884
tri 20964 47602 21246 47884 sw
tri 21246 47602 21528 47884 ne
rect 21528 47780 25297 47884
tri 25297 47780 25594 48077 sw
tri 25594 47780 25891 48077 ne
rect 25891 47802 27560 48077
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48090 29540 48091
tri 29540 48090 29830 48380 sw
tri 29830 48090 30120 48380 ne
rect 30120 48314 33846 48380
tri 33846 48314 34140 48608 sw
tri 34140 48314 34434 48608 ne
rect 34434 48448 38256 48608
tri 38256 48448 38544 48736 sw
tri 38544 48448 38832 48736 ne
rect 38832 48538 42689 48736
tri 42689 48538 42986 48835 sw
tri 42986 48538 43283 48835 ne
rect 43283 48627 47145 48835
tri 47145 48627 47438 48920 sw
tri 47438 48627 47731 48920 ne
rect 47731 48832 49418 48920
tri 49418 48832 49506 48920 sw
tri 49710 48832 49798 48920 ne
rect 49798 48845 51478 48920
tri 51478 48845 51765 49132 sw
tri 51765 48845 52052 49132 ne
rect 52052 49005 55834 49132
tri 55834 49005 56145 49316 sw
tri 56145 49005 56456 49316 ne
rect 56456 49200 60225 49316
tri 60225 49200 60510 49485 sw
tri 60510 49200 60795 49485 ne
rect 60795 49200 71000 49485
rect 56456 49005 60510 49200
rect 52052 48845 56145 49005
rect 49798 48832 51765 48845
rect 47731 48627 49506 48832
rect 43283 48538 47438 48627
rect 38832 48448 42986 48538
rect 34434 48416 38544 48448
tri 38544 48416 38576 48448 sw
tri 38832 48416 38864 48448 ne
rect 38864 48416 42986 48448
rect 34434 48314 38576 48416
rect 30120 48090 34140 48314
rect 28138 48020 29830 48090
tri 29830 48020 29900 48090 sw
tri 30120 48020 30190 48090 ne
rect 30190 48020 34140 48090
tri 34140 48020 34434 48314 sw
tri 34434 48020 34728 48314 ne
rect 34728 48128 38576 48314
tri 38576 48128 38864 48416 sw
tri 38864 48128 39152 48416 ne
rect 39152 48241 42986 48416
tri 42986 48241 43283 48538 sw
tri 43283 48241 43580 48538 ne
rect 43580 48334 47438 48538
tri 47438 48334 47731 48627 sw
tri 47731 48334 48024 48627 ne
rect 48024 48540 49506 48627
tri 49506 48540 49798 48832 sw
tri 49798 48540 50090 48832 ne
rect 50090 48827 51765 48832
tri 51765 48827 51783 48845 sw
tri 52052 48827 52070 48845 ne
rect 52070 48827 56145 48845
rect 50090 48540 51783 48827
tri 51783 48540 52070 48827 sw
tri 52070 48540 52357 48827 ne
rect 52357 48694 56145 48827
tri 56145 48694 56456 49005 sw
tri 56456 48694 56767 49005 ne
rect 56767 49000 60510 49005
tri 60510 49000 60710 49200 sw
rect 56767 48694 71000 49000
rect 52357 48608 56456 48694
tri 56456 48608 56542 48694 sw
tri 56767 48608 56853 48694 ne
rect 56853 48608 71000 48694
rect 52357 48540 56542 48608
rect 48024 48334 49798 48540
rect 43580 48241 47731 48334
rect 39152 48128 43283 48241
rect 34728 48020 38864 48128
rect 28138 47802 29900 48020
rect 25891 47780 27849 47802
rect 21528 47671 25594 47780
tri 25594 47671 25703 47780 sw
tri 25891 47671 26000 47780 ne
rect 26000 47671 27849 47780
rect 21528 47602 25703 47671
rect 17200 47404 21246 47602
tri 17200 47312 17292 47404 ne
rect 17292 47320 21246 47404
tri 21246 47320 21528 47602 sw
tri 21528 47320 21810 47602 ne
rect 21810 47374 25703 47602
tri 25703 47374 26000 47671 sw
tri 26000 47374 26297 47671 ne
rect 26297 47513 27849 47671
tri 27849 47513 28138 47802 sw
tri 28138 47513 28427 47802 ne
rect 28427 47730 29900 47802
tri 29900 47730 30190 48020 sw
tri 30190 47730 30480 48020 ne
rect 30480 47730 34434 48020
rect 28427 47513 30190 47730
rect 26297 47374 28138 47513
rect 21810 47320 26000 47374
rect 17292 47312 21528 47320
tri 17000 47112 17200 47312 sw
tri 17292 47112 17492 47312 ne
rect 17492 47274 21528 47312
tri 21528 47274 21574 47320 sw
tri 21810 47274 21856 47320 ne
rect 21856 47274 26000 47320
rect 17492 47112 21574 47274
rect 14000 46908 17200 47112
tri 17200 46908 17404 47112 sw
tri 17492 46908 17696 47112 ne
rect 17696 46992 21574 47112
tri 21574 46992 21856 47274 sw
tri 21856 46992 22138 47274 ne
rect 22138 47077 26000 47274
tri 26000 47077 26297 47374 sw
tri 26297 47077 26594 47374 ne
rect 26594 47358 28138 47374
tri 28138 47358 28293 47513 sw
tri 28427 47358 28582 47513 ne
rect 28582 47440 30190 47513
tri 30190 47440 30480 47730 sw
tri 30480 47440 30770 47730 ne
rect 30770 47726 34434 47730
tri 34434 47726 34728 48020 sw
tri 34728 47726 35022 48020 ne
rect 35022 47840 38864 48020
tri 38864 47840 39152 48128 sw
tri 39152 47840 39440 48128 ne
rect 39440 47944 43283 48128
tri 43283 47944 43580 48241 sw
tri 43580 47944 43877 48241 ne
rect 43877 48041 47731 48241
tri 47731 48041 48024 48334 sw
tri 48024 48041 48317 48334 ne
rect 48317 48248 49798 48334
tri 49798 48248 50090 48540 sw
tri 50090 48248 50382 48540 ne
rect 50382 48253 52070 48540
tri 52070 48253 52357 48540 sw
tri 52357 48253 52644 48540 ne
rect 52644 48297 56542 48540
tri 56542 48297 56853 48608 sw
tri 56853 48297 57164 48608 ne
rect 57164 48297 71000 48608
rect 52644 48253 56853 48297
rect 50382 48248 52357 48253
rect 48317 48041 50090 48248
rect 43877 47944 48024 48041
rect 39440 47840 43580 47944
rect 35022 47726 39152 47840
rect 30770 47564 34728 47726
tri 34728 47564 34890 47726 sw
tri 35022 47564 35184 47726 ne
rect 35184 47564 39152 47726
rect 30770 47440 34890 47564
rect 28582 47358 30480 47440
rect 26594 47077 28293 47358
rect 22138 46992 26297 47077
rect 17696 46908 21856 46992
rect 14000 46616 17404 46908
tri 17404 46616 17696 46908 sw
tri 17696 46616 17988 46908 ne
rect 17988 46710 21856 46908
tri 21856 46710 22138 46992 sw
tri 22138 46710 22420 46992 ne
rect 22420 46780 26297 46992
tri 26297 46780 26594 47077 sw
tri 26594 46780 26891 47077 ne
rect 26891 47069 28293 47077
tri 28293 47069 28582 47358 sw
tri 28582 47069 28871 47358 ne
rect 28871 47266 30480 47358
tri 30480 47266 30654 47440 sw
tri 30770 47266 30944 47440 ne
rect 30944 47270 34890 47440
tri 34890 47270 35184 47564 sw
tri 35184 47270 35478 47564 ne
rect 35478 47552 39152 47564
tri 39152 47552 39440 47840 sw
tri 39440 47552 39728 47840 ne
rect 39728 47647 43580 47840
tri 43580 47647 43877 47944 sw
tri 43877 47647 44174 47944 ne
rect 44174 47819 48024 47944
tri 48024 47819 48246 48041 sw
tri 48317 47819 48539 48041 ne
rect 48539 47956 50090 48041
tri 50090 47956 50382 48248 sw
tri 50382 47956 50674 48248 ne
rect 50674 47966 52357 48248
tri 52357 47966 52644 48253 sw
tri 52644 47966 52931 48253 ne
rect 52931 47986 56853 48253
tri 56853 47986 57164 48297 sw
tri 57164 47986 57475 48297 ne
rect 57475 47986 71000 48297
rect 52931 47966 57164 47986
rect 50674 47956 52644 47966
rect 48539 47819 50382 47956
rect 44174 47647 48246 47819
rect 39728 47552 43877 47647
rect 35478 47270 39440 47552
rect 30944 47266 35184 47270
rect 28871 47069 30654 47266
rect 26891 46780 28582 47069
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 46976 30654 47069
tri 30654 46976 30944 47266 sw
tri 30944 46976 31234 47266 ne
rect 31234 46976 35184 47266
tri 35184 46976 35478 47270 sw
tri 35478 46976 35772 47270 ne
rect 35772 47264 39440 47270
tri 39440 47264 39728 47552 sw
tri 39728 47264 40016 47552 ne
rect 40016 47417 43877 47552
tri 43877 47417 44107 47647 sw
tri 44174 47417 44404 47647 ne
rect 44404 47526 48246 47647
tri 48246 47526 48539 47819 sw
tri 48539 47526 48832 47819 ne
rect 48832 47664 50382 47819
tri 50382 47664 50674 47956 sw
tri 50674 47664 50966 47956 ne
rect 50966 47679 52644 47956
tri 52644 47679 52931 47966 sw
tri 52931 47679 53218 47966 ne
rect 53218 47679 57164 47966
rect 50966 47664 52931 47679
rect 48832 47526 50674 47664
rect 44404 47417 48539 47526
rect 40016 47264 44107 47417
rect 35772 46976 39728 47264
tri 39728 46976 40016 47264 sw
tri 40016 46976 40304 47264 ne
rect 40304 47120 44107 47264
tri 44107 47120 44404 47417 sw
tri 44404 47120 44701 47417 ne
rect 44701 47233 48539 47417
tri 48539 47233 48832 47526 sw
tri 48832 47233 49125 47526 ne
rect 49125 47524 50674 47526
tri 50674 47524 50814 47664 sw
tri 50966 47524 51106 47664 ne
rect 51106 47627 52931 47664
tri 52931 47627 52983 47679 sw
tri 53218 47627 53270 47679 ne
rect 53270 47675 57164 47679
tri 57164 47675 57475 47986 sw
tri 57475 47675 57786 47986 ne
rect 57786 47675 71000 47986
rect 53270 47627 57475 47675
rect 51106 47524 52983 47627
rect 49125 47233 50814 47524
rect 44701 47120 48832 47233
rect 40304 46976 44404 47120
rect 29160 46780 30944 46976
rect 22420 46710 26594 46780
rect 17988 46616 22138 46710
rect 14000 46324 17696 46616
tri 17696 46324 17988 46616 sw
tri 17988 46324 18280 46616 ne
rect 18280 46428 22138 46616
tri 22138 46428 22420 46710 sw
tri 22420 46428 22702 46710 ne
rect 22702 46483 26594 46710
tri 26594 46483 26891 46780 sw
tri 26891 46483 27188 46780 ne
rect 27188 46689 28871 46780
tri 28871 46689 28962 46780 sw
tri 29160 46689 29251 46780 ne
rect 29251 46690 30944 46780
tri 30944 46690 31230 46976 sw
tri 31234 46690 31520 46976 ne
rect 31520 46690 35478 46976
rect 29251 46689 31230 46690
rect 27188 46483 28962 46689
rect 22702 46428 26891 46483
rect 18280 46324 22420 46428
rect 14000 46068 17988 46324
tri 14000 42497 17571 46068 ne
rect 17571 46032 17988 46068
tri 17988 46032 18280 46324 sw
tri 18280 46032 18572 46324 ne
rect 18572 46146 22420 46324
tri 22420 46146 22702 46428 sw
tri 22702 46146 22984 46428 ne
rect 22984 46186 26891 46428
tri 26891 46186 27188 46483 sw
tri 27188 46186 27485 46483 ne
rect 27485 46400 28962 46483
tri 28962 46400 29251 46689 sw
tri 29251 46400 29540 46689 ne
rect 29540 46400 31230 46689
tri 31230 46400 31520 46690 sw
tri 31520 46400 31810 46690 ne
rect 31810 46682 35478 46690
tri 35478 46682 35772 46976 sw
tri 35772 46682 36066 46976 ne
rect 36066 46688 40016 46976
tri 40016 46688 40304 46976 sw
tri 40304 46688 40592 46976 ne
rect 40592 46823 44404 46976
tri 44404 46823 44701 47120 sw
tri 44701 46823 44998 47120 ne
rect 44998 46940 48832 47120
tri 48832 46940 49125 47233 sw
tri 49125 46940 49418 47233 ne
rect 49418 47232 50814 47233
tri 50814 47232 51106 47524 sw
tri 51106 47232 51398 47524 ne
rect 51398 47340 52983 47524
tri 52983 47340 53270 47627 sw
tri 53270 47340 53557 47627 ne
rect 53557 47364 57475 47627
tri 57475 47364 57786 47675 sw
tri 57786 47364 58097 47675 ne
rect 58097 47364 71000 47675
rect 53557 47340 57786 47364
rect 51398 47232 53270 47340
rect 49418 46940 51106 47232
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47053 53270 47232
tri 53270 47053 53557 47340 sw
tri 53557 47053 53844 47340 ne
rect 53844 47053 57786 47340
tri 57786 47053 58097 47364 sw
tri 58097 47053 58408 47364 ne
rect 58408 47053 71000 47364
rect 51690 46940 53557 47053
rect 44998 46823 49125 46940
rect 40592 46688 44701 46823
rect 36066 46682 40304 46688
rect 31810 46400 35772 46682
rect 27485 46186 29251 46400
rect 22984 46146 27188 46186
rect 18572 46032 22702 46146
rect 17571 45740 18280 46032
tri 18280 45740 18572 46032 sw
tri 18572 45740 18864 46032 ne
rect 18864 45864 22702 46032
tri 22702 45864 22984 46146 sw
tri 22984 45864 23266 46146 ne
rect 23266 45889 27188 46146
tri 27188 45889 27485 46186 sw
tri 27485 45889 27782 46186 ne
rect 27782 46111 29251 46186
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46111 31520 46400
rect 27782 45889 29540 46111
rect 23266 45864 27485 45889
rect 18864 45740 22984 45864
rect 17571 45448 18572 45740
tri 18572 45448 18864 45740 sw
tri 18864 45448 19156 45740 ne
rect 19156 45582 22984 45740
tri 22984 45582 23266 45864 sw
tri 23266 45582 23548 45864 ne
rect 23548 45691 27485 45864
tri 27485 45691 27683 45889 sw
tri 27782 45691 27980 45889 ne
rect 27980 45822 29540 45889
tri 29540 45822 29829 46111 sw
tri 29829 45822 30118 46111 ne
rect 30118 46110 31520 46111
tri 31520 46110 31810 46400 sw
tri 31810 46110 32100 46400 ne
rect 32100 46388 35772 46400
tri 35772 46388 36066 46682 sw
tri 36066 46388 36360 46682 ne
rect 36360 46508 40304 46682
tri 40304 46508 40484 46688 sw
tri 40592 46508 40772 46688 ne
rect 40772 46526 44701 46688
tri 44701 46526 44998 46823 sw
tri 44998 46526 45295 46823 ne
rect 45295 46647 49125 46823
tri 49125 46647 49418 46940 sw
tri 49418 46647 49711 46940 ne
rect 49711 46852 51398 46940
tri 51398 46852 51486 46940 sw
tri 51690 46852 51778 46940 ne
rect 51778 46852 53557 46940
rect 49711 46647 51486 46852
rect 45295 46526 49418 46647
rect 40772 46508 44998 46526
rect 36360 46388 40484 46508
rect 32100 46110 36066 46388
rect 30118 45864 31810 46110
tri 31810 45864 32056 46110 sw
tri 32100 45864 32346 46110 ne
rect 32346 46094 36066 46110
tri 36066 46094 36360 46388 sw
tri 36360 46094 36654 46388 ne
rect 36654 46220 40484 46388
tri 40484 46220 40772 46508 sw
tri 40772 46220 41060 46508 ne
rect 41060 46229 44998 46508
tri 44998 46229 45295 46526 sw
tri 45295 46229 45592 46526 ne
rect 45592 46354 49418 46526
tri 49418 46354 49711 46647 sw
tri 49711 46354 50004 46647 ne
rect 50004 46560 51486 46647
tri 51486 46560 51778 46852 sw
tri 51778 46560 52070 46852 ne
rect 52070 46847 53557 46852
tri 53557 46847 53763 47053 sw
tri 53844 46847 54050 47053 ne
rect 54050 46847 58097 47053
rect 52070 46560 53763 46847
tri 53763 46560 54050 46847 sw
tri 54050 46560 54337 46847 ne
rect 54337 46742 58097 46847
tri 58097 46742 58408 47053 sw
tri 58408 46742 58719 47053 ne
rect 58719 46742 71000 47053
rect 54337 46622 58408 46742
tri 58408 46622 58528 46742 sw
tri 58719 46622 58839 46742 ne
rect 58839 46622 71000 46742
rect 54337 46560 58528 46622
rect 50004 46354 51778 46560
rect 45592 46229 49711 46354
rect 41060 46220 45295 46229
rect 36654 46094 40772 46220
rect 32346 45864 36360 46094
rect 30118 45822 32056 45864
rect 27980 45691 29829 45822
rect 23548 45582 27683 45691
rect 19156 45448 23266 45582
rect 17571 45168 18864 45448
tri 18864 45168 19144 45448 sw
tri 19156 45168 19436 45448 ne
rect 19436 45300 23266 45448
tri 23266 45300 23548 45582 sw
tri 23548 45300 23830 45582 ne
rect 23830 45394 27683 45582
tri 27683 45394 27980 45691 sw
tri 27980 45394 28277 45691 ne
rect 28277 45533 29829 45691
tri 29829 45533 30118 45822 sw
tri 30118 45533 30407 45822 ne
rect 30407 45574 32056 45822
tri 32056 45574 32346 45864 sw
tri 32346 45574 32636 45864 ne
rect 32636 45800 36360 45864
tri 36360 45800 36654 46094 sw
tri 36654 45800 36948 46094 ne
rect 36948 45932 40772 46094
tri 40772 45932 41060 46220 sw
tri 41060 45932 41348 46220 ne
rect 41348 45932 45295 46220
tri 45295 45932 45592 46229 sw
tri 45592 45932 45889 46229 ne
rect 45889 46061 49711 46229
tri 49711 46061 50004 46354 sw
tri 50004 46061 50297 46354 ne
rect 50297 46268 51778 46354
tri 51778 46268 52070 46560 sw
tri 52070 46268 52362 46560 ne
rect 52362 46273 54050 46560
tri 54050 46273 54337 46560 sw
tri 54337 46273 54624 46560 ne
rect 54624 46311 58528 46560
tri 58528 46311 58839 46622 sw
tri 58839 46311 59150 46622 ne
rect 59150 46311 71000 46622
rect 54624 46273 58839 46311
rect 52362 46268 54337 46273
rect 50297 46061 52070 46268
rect 45889 45932 50004 46061
rect 36948 45800 41060 45932
rect 32636 45574 36654 45800
rect 30407 45533 32346 45574
rect 28277 45394 30118 45533
rect 23830 45300 27980 45394
rect 19436 45168 23548 45300
rect 17571 44876 19144 45168
tri 19144 44876 19436 45168 sw
tri 19436 44876 19728 45168 ne
rect 19728 45018 23548 45168
tri 23548 45018 23830 45300 sw
tri 23830 45018 24112 45300 ne
rect 24112 45097 27980 45300
tri 27980 45097 28277 45394 sw
tri 28277 45097 28574 45394 ne
rect 28574 45378 30118 45394
tri 30118 45378 30273 45533 sw
tri 30407 45378 30562 45533 ne
rect 30562 45378 32346 45533
rect 28574 45097 30273 45378
rect 24112 45018 28277 45097
rect 19728 44876 23830 45018
rect 17571 44584 19436 44876
tri 19436 44584 19728 44876 sw
tri 19728 44584 20020 44876 ne
rect 20020 44736 23830 44876
tri 23830 44736 24112 45018 sw
tri 24112 44736 24394 45018 ne
rect 24394 44800 28277 45018
tri 28277 44800 28574 45097 sw
tri 28574 44800 28871 45097 ne
rect 28871 45089 30273 45097
tri 30273 45089 30562 45378 sw
tri 30562 45089 30851 45378 ne
rect 30851 45284 32346 45378
tri 32346 45284 32636 45574 sw
tri 32636 45284 32926 45574 ne
rect 32926 45506 36654 45574
tri 36654 45506 36948 45800 sw
tri 36948 45506 37242 45800 ne
rect 37242 45644 41060 45800
tri 41060 45644 41348 45932 sw
tri 41348 45644 41636 45932 ne
rect 41636 45644 45592 45932
rect 37242 45506 41348 45644
rect 32926 45284 36948 45506
rect 30851 45089 32636 45284
rect 28871 44800 30562 45089
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 45000 32636 45089
tri 32636 45000 32920 45284 sw
tri 32926 45000 33210 45284 ne
rect 33210 45246 36948 45284
tri 36948 45246 37208 45506 sw
tri 37242 45246 37502 45506 ne
rect 37502 45356 41348 45506
tri 41348 45356 41636 45644 sw
tri 41636 45356 41924 45644 ne
rect 41924 45635 45592 45644
tri 45592 45635 45889 45932 sw
tri 45889 45635 46186 45932 ne
rect 46186 45839 50004 45932
tri 50004 45839 50226 46061 sw
tri 50297 45839 50519 46061 ne
rect 50519 45976 52070 46061
tri 52070 45976 52362 46268 sw
tri 52362 45976 52654 46268 ne
rect 52654 46000 54337 46268
tri 54337 46000 54610 46273 sw
tri 54624 46000 54897 46273 ne
rect 54897 46000 58839 46273
tri 58839 46000 59150 46311 sw
tri 59150 46000 59461 46311 ne
rect 59461 46000 71000 46311
rect 52654 45976 54610 46000
rect 50519 45839 52362 45976
rect 46186 45635 50226 45839
rect 41924 45482 45889 45635
tri 45889 45482 46042 45635 sw
tri 46186 45482 46339 45635 ne
rect 46339 45546 50226 45635
tri 50226 45546 50519 45839 sw
tri 50519 45546 50812 45839 ne
rect 50812 45684 52362 45839
tri 52362 45684 52654 45976 sw
tri 52654 45684 52946 45976 ne
rect 52946 45713 54610 45976
tri 54610 45713 54897 46000 sw
tri 54897 45713 55184 46000 ne
rect 55184 45799 59150 46000
tri 59150 45799 59351 46000 sw
rect 55184 45739 71000 45799
rect 55184 45713 70613 45739
rect 52946 45684 54897 45713
rect 50812 45546 52654 45684
rect 46339 45482 50519 45546
rect 41924 45356 46042 45482
rect 37502 45246 41636 45356
rect 33210 45000 37208 45246
rect 31140 44800 32920 45000
rect 24394 44736 28574 44800
rect 20020 44584 24112 44736
rect 17571 44292 19728 44584
tri 19728 44292 20020 44584 sw
tri 20020 44292 20312 44584 ne
rect 20312 44454 24112 44584
tri 24112 44454 24394 44736 sw
tri 24394 44454 24676 44736 ne
rect 24676 44503 28574 44736
tri 28574 44503 28871 44800 sw
tri 28871 44503 29168 44800 ne
rect 29168 44709 30851 44800
tri 30851 44709 30942 44800 sw
tri 31140 44709 31231 44800 ne
rect 31231 44710 32920 44800
tri 32920 44710 33210 45000 sw
tri 33210 44710 33500 45000 ne
rect 33500 44952 37208 45000
tri 37208 44952 37502 45246 sw
tri 37502 44952 37796 45246 ne
rect 37796 45068 41636 45246
tri 41636 45068 41924 45356 sw
tri 41924 45068 42212 45356 ne
rect 42212 45185 46042 45356
tri 46042 45185 46339 45482 sw
tri 46339 45185 46636 45482 ne
rect 46636 45253 50519 45482
tri 50519 45253 50812 45546 sw
tri 50812 45253 51105 45546 ne
rect 51105 45472 52654 45546
tri 52654 45472 52866 45684 sw
tri 52946 45472 53158 45684 ne
rect 53158 45472 54897 45684
rect 51105 45253 52866 45472
rect 46636 45185 50812 45253
rect 42212 45068 46339 45185
rect 37796 44952 41924 45068
rect 33500 44710 37502 44952
rect 31231 44709 33210 44710
rect 29168 44503 30942 44709
rect 24676 44454 28871 44503
rect 20312 44292 24394 44454
rect 17571 44000 20020 44292
tri 20020 44000 20312 44292 sw
tri 20312 44000 20604 44292 ne
rect 20604 44172 24394 44292
tri 24394 44172 24676 44454 sw
tri 24676 44172 24958 44454 ne
rect 24958 44206 28871 44454
tri 28871 44206 29168 44503 sw
tri 29168 44206 29465 44503 ne
rect 29465 44420 30942 44503
tri 30942 44420 31231 44709 sw
tri 31231 44420 31520 44709 ne
rect 31520 44420 33210 44709
tri 33210 44420 33500 44710 sw
tri 33500 44420 33790 44710 ne
rect 33790 44658 37502 44710
tri 37502 44658 37796 44952 sw
tri 37796 44658 38090 44952 ne
rect 38090 44780 41924 44952
tri 41924 44780 42212 45068 sw
tri 42212 44780 42500 45068 ne
rect 42500 44888 46339 45068
tri 46339 44888 46636 45185 sw
tri 46636 44888 46933 45185 ne
rect 46933 44960 50812 45185
tri 50812 44960 51105 45253 sw
tri 51105 44960 51398 45253 ne
rect 51398 45180 52866 45253
tri 52866 45180 53158 45472 sw
tri 53158 45180 53450 45472 ne
rect 53450 45426 54897 45472
tri 54897 45426 55184 45713 sw
tri 55184 45426 55471 45713 ne
rect 55471 45426 70613 45713
rect 53450 45180 55184 45426
rect 51398 44960 53158 45180
rect 46933 44888 51105 44960
rect 42500 44780 46636 44888
rect 38090 44658 42212 44780
rect 33790 44420 37796 44658
rect 29465 44206 31231 44420
rect 24958 44172 29168 44206
rect 20604 44000 24676 44172
rect 17571 43708 20312 44000
tri 20312 43708 20604 44000 sw
tri 20604 43708 20896 44000 ne
rect 20896 43917 24676 44000
tri 24676 43917 24931 44172 sw
tri 24958 43917 25213 44172 ne
rect 25213 43917 29168 44172
rect 20896 43708 24931 43917
rect 17571 43416 20604 43708
tri 20604 43416 20896 43708 sw
tri 20896 43416 21188 43708 ne
rect 21188 43635 24931 43708
tri 24931 43635 25213 43917 sw
tri 25213 43635 25495 43917 ne
rect 25495 43909 29168 43917
tri 29168 43909 29465 44206 sw
tri 29465 43909 29762 44206 ne
rect 29762 44131 31231 44206
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44131 33500 44420
rect 29762 43909 31520 44131
rect 25495 43711 29465 43909
tri 29465 43711 29663 43909 sw
tri 29762 43711 29960 43909 ne
rect 29960 43842 31520 43909
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44130 33500 44131
tri 33500 44130 33790 44420 sw
tri 33790 44130 34080 44420 ne
rect 34080 44364 37796 44420
tri 37796 44364 38090 44658 sw
tri 38090 44364 38384 44658 ne
rect 38384 44492 42212 44658
tri 42212 44492 42500 44780 sw
tri 42500 44492 42788 44780 ne
rect 42788 44591 46636 44780
tri 46636 44591 46933 44888 sw
tri 46933 44591 47230 44888 ne
rect 47230 44667 51105 44888
tri 51105 44667 51398 44960 sw
tri 51398 44667 51691 44960 ne
rect 51691 44888 53158 44960
tri 53158 44888 53450 45180 sw
tri 53450 44888 53742 45180 ne
rect 53742 45175 55184 45180
tri 55184 45175 55435 45426 sw
tri 55471 45175 55722 45426 ne
rect 55722 45175 70613 45426
rect 53742 44888 55435 45175
tri 55435 44888 55722 45175 sw
tri 55722 44888 56009 45175 ne
rect 56009 44888 70613 45175
rect 51691 44872 53450 44888
tri 53450 44872 53466 44888 sw
tri 53742 44872 53758 44888 ne
rect 53758 44872 55722 44888
rect 51691 44667 53466 44872
rect 47230 44591 51398 44667
rect 42788 44492 46933 44591
rect 38384 44364 42500 44492
rect 34080 44130 38090 44364
rect 32098 44066 33790 44130
tri 33790 44066 33854 44130 sw
tri 34080 44066 34144 44130 ne
rect 34144 44070 38090 44130
tri 38090 44070 38384 44364 sw
tri 38384 44070 38678 44364 ne
rect 38678 44204 42500 44364
tri 42500 44204 42788 44492 sw
tri 42788 44204 43076 44492 ne
rect 43076 44294 46933 44492
tri 46933 44294 47230 44591 sw
tri 47230 44294 47527 44591 ne
rect 47527 44374 51398 44591
tri 51398 44374 51691 44667 sw
tri 51691 44374 51984 44667 ne
rect 51984 44580 53466 44667
tri 53466 44580 53758 44872 sw
tri 53758 44580 54050 44872 ne
rect 54050 44867 55722 44872
tri 55722 44867 55743 44888 sw
tri 56009 44867 56030 44888 ne
rect 56030 44867 70613 44888
rect 54050 44580 55743 44867
tri 55743 44580 56030 44867 sw
tri 56030 44580 56317 44867 ne
rect 56317 44580 70613 44867
rect 51984 44374 53758 44580
rect 47527 44294 51691 44374
rect 43076 44204 47230 44294
rect 38678 44172 42788 44204
tri 42788 44172 42820 44204 sw
tri 43076 44172 43108 44204 ne
rect 43108 44172 47230 44204
rect 38678 44070 42820 44172
rect 34144 44066 38384 44070
rect 32098 43842 33854 44066
rect 29960 43711 31809 43842
rect 25495 43635 29663 43711
rect 21188 43416 25213 43635
rect 17571 43248 20896 43416
tri 20896 43248 21064 43416 sw
tri 21188 43248 21356 43416 ne
rect 21356 43353 25213 43416
tri 25213 43353 25495 43635 sw
tri 25495 43353 25777 43635 ne
rect 25777 43414 29663 43635
tri 29663 43414 29960 43711 sw
tri 29960 43414 30257 43711 ne
rect 30257 43553 31809 43711
tri 31809 43553 32098 43842 sw
tri 32098 43553 32387 43842 ne
rect 32387 43776 33854 43842
tri 33854 43776 34144 44066 sw
tri 34144 43776 34434 44066 ne
rect 34434 43776 38384 44066
tri 38384 43776 38678 44070 sw
tri 38678 43776 38972 44070 ne
rect 38972 43884 42820 44070
tri 42820 43884 43108 44172 sw
tri 43108 43884 43396 44172 ne
rect 43396 43997 47230 44172
tri 47230 43997 47527 44294 sw
tri 47527 43997 47824 44294 ne
rect 47824 44081 51691 44294
tri 51691 44081 51984 44374 sw
tri 51984 44081 52277 44374 ne
rect 52277 44288 53758 44374
tri 53758 44288 54050 44580 sw
tri 54050 44288 54342 44580 ne
rect 54342 44293 56030 44580
tri 56030 44293 56317 44580 sw
tri 56317 44293 56604 44580 ne
rect 56604 44293 70613 44580
rect 54342 44288 56317 44293
rect 52277 44081 54050 44288
rect 47824 43997 51984 44081
rect 43396 43884 47527 43997
rect 38972 43776 43108 43884
rect 32387 43553 34144 43776
rect 30257 43414 32098 43553
rect 25777 43353 29960 43414
rect 21356 43248 25495 43353
rect 17571 42956 21064 43248
tri 21064 42956 21356 43248 sw
tri 21356 42956 21648 43248 ne
rect 21648 43071 25495 43248
tri 25495 43071 25777 43353 sw
tri 25777 43071 26059 43353 ne
rect 26059 43117 29960 43353
tri 29960 43117 30257 43414 sw
tri 30257 43117 30554 43414 ne
rect 30554 43398 32098 43414
tri 32098 43398 32253 43553 sw
tri 32387 43398 32542 43553 ne
rect 32542 43486 34144 43553
tri 34144 43486 34434 43776 sw
tri 34434 43486 34724 43776 ne
rect 34724 43486 38678 43776
rect 32542 43398 34434 43486
rect 30554 43117 32253 43398
rect 26059 43071 30257 43117
rect 21648 42956 25777 43071
rect 17571 42664 21356 42956
tri 21356 42664 21648 42956 sw
tri 21648 42664 21940 42956 ne
rect 21940 42789 25777 42956
tri 25777 42789 26059 43071 sw
tri 26059 42789 26341 43071 ne
rect 26341 42820 30257 43071
tri 30257 42820 30554 43117 sw
tri 30554 42820 30851 43117 ne
rect 30851 43109 32253 43117
tri 32253 43109 32542 43398 sw
tri 32542 43109 32831 43398 ne
rect 32831 43196 34434 43398
tri 34434 43196 34724 43486 sw
tri 34724 43196 35014 43486 ne
rect 35014 43482 38678 43486
tri 38678 43482 38972 43776 sw
tri 38972 43482 39266 43776 ne
rect 39266 43596 43108 43776
tri 43108 43596 43396 43884 sw
tri 43396 43596 43684 43884 ne
rect 43684 43700 47527 43884
tri 47527 43700 47824 43997 sw
tri 47824 43700 48121 43997 ne
rect 48121 43859 51984 43997
tri 51984 43859 52206 44081 sw
tri 52277 43859 52499 44081 ne
rect 52499 43996 54050 44081
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44006 56317 44288
tri 56317 44006 56604 44293 sw
tri 56604 44006 56891 44293 ne
rect 56891 44006 70613 44293
rect 54634 43996 56604 44006
rect 52499 43859 54342 43996
rect 48121 43700 52206 43859
rect 43684 43596 47824 43700
rect 39266 43482 43396 43596
rect 35014 43320 38972 43482
tri 38972 43320 39134 43482 sw
tri 39266 43320 39428 43482 ne
rect 39428 43320 43396 43482
rect 35014 43196 39134 43320
rect 32831 43109 34724 43196
rect 30851 42820 32542 43109
tri 32542 42820 32831 43109 sw
tri 32831 42820 33120 43109 ne
rect 33120 43020 34724 43109
tri 34724 43020 34900 43196 sw
tri 35014 43020 35190 43196 ne
rect 35190 43026 39134 43196
tri 39134 43026 39428 43320 sw
tri 39428 43026 39722 43320 ne
rect 39722 43308 43396 43320
tri 43396 43308 43684 43596 sw
tri 43684 43308 43972 43596 ne
rect 43972 43403 47824 43596
tri 47824 43403 48121 43700 sw
tri 48121 43403 48418 43700 ne
rect 48418 43566 52206 43700
tri 52206 43566 52499 43859 sw
tri 52499 43566 52792 43859 ne
rect 52792 43704 54342 43859
tri 54342 43704 54634 43996 sw
tri 54634 43704 54926 43996 ne
rect 54926 43719 56604 43996
tri 56604 43719 56891 44006 sw
tri 56891 43719 57178 44006 ne
rect 57178 43719 70613 44006
rect 54926 43704 56891 43719
rect 52792 43676 54634 43704
tri 54634 43676 54662 43704 sw
tri 54926 43676 54954 43704 ne
rect 54954 43676 56891 43704
rect 52792 43566 54662 43676
rect 48418 43403 52499 43566
rect 43972 43308 48121 43403
rect 39722 43026 43684 43308
rect 35190 43020 39428 43026
rect 33120 42820 34900 43020
rect 26341 42789 30554 42820
rect 21940 42664 26059 42789
rect 17571 42497 21648 42664
tri 17571 38420 21648 42497 ne
tri 21648 42372 21940 42664 sw
tri 21940 42372 22232 42664 ne
rect 22232 42507 26059 42664
tri 26059 42507 26341 42789 sw
tri 26341 42507 26623 42789 ne
rect 26623 42523 30554 42789
tri 30554 42523 30851 42820 sw
tri 30851 42523 31148 42820 ne
rect 31148 42729 32831 42820
tri 32831 42729 32922 42820 sw
tri 33120 42729 33211 42820 ne
rect 33211 42730 34900 42820
tri 34900 42730 35190 43020 sw
tri 35190 42730 35480 43020 ne
rect 35480 42732 39428 43020
tri 39428 42732 39722 43026 sw
tri 39722 42732 40016 43026 ne
rect 40016 43020 43684 43026
tri 43684 43020 43972 43308 sw
tri 43972 43020 44260 43308 ne
rect 44260 43173 48121 43308
tri 48121 43173 48351 43403 sw
tri 48418 43173 48648 43403 ne
rect 48648 43273 52499 43403
tri 52499 43273 52792 43566 sw
tri 52792 43273 53085 43566 ne
rect 53085 43384 54662 43566
tri 54662 43384 54954 43676 sw
tri 54954 43384 55246 43676 ne
rect 55246 43461 56891 43676
tri 56891 43461 57149 43719 sw
tri 57178 43461 57436 43719 ne
rect 57436 43461 70613 43719
rect 55246 43384 57149 43461
rect 53085 43273 54954 43384
rect 48648 43173 52792 43273
rect 44260 43020 48351 43173
rect 40016 42732 43972 43020
tri 43972 42732 44260 43020 sw
tri 44260 42732 44548 43020 ne
rect 44548 42876 48351 43020
tri 48351 42876 48648 43173 sw
tri 48648 42876 48945 43173 ne
rect 48945 42980 52792 43173
tri 52792 42980 53085 43273 sw
tri 53085 42980 53378 43273 ne
rect 53378 43092 54954 43273
tri 54954 43092 55246 43384 sw
tri 55246 43092 55538 43384 ne
rect 55538 43174 57149 43384
tri 57149 43174 57436 43461 sw
tri 57436 43174 57723 43461 ne
rect 57723 43174 70613 43461
rect 55538 43092 57436 43174
rect 53378 42980 55246 43092
rect 48945 42876 53085 42980
rect 44548 42732 48648 42876
rect 35480 42730 39722 42732
rect 33211 42729 35190 42730
rect 31148 42523 32922 42729
rect 26623 42507 30851 42523
rect 22232 42372 26341 42507
rect 21648 42080 21940 42372
tri 21940 42080 22232 42372 sw
tri 22232 42080 22524 42372 ne
rect 22524 42225 26341 42372
tri 26341 42225 26623 42507 sw
tri 26623 42225 26905 42507 ne
rect 26905 42226 30851 42507
tri 30851 42226 31148 42523 sw
tri 31148 42226 31445 42523 ne
rect 31445 42440 32922 42523
tri 32922 42440 33211 42729 sw
tri 33211 42440 33500 42729 ne
rect 33500 42440 35190 42729
tri 35190 42440 35480 42730 sw
tri 35480 42440 35770 42730 ne
rect 35770 42440 39722 42730
rect 31445 42226 33211 42440
rect 26905 42225 31148 42226
rect 22524 42184 26623 42225
tri 26623 42184 26664 42225 sw
tri 26905 42184 26946 42225 ne
rect 26946 42184 31148 42225
rect 22524 42080 26664 42184
rect 21648 41788 22232 42080
tri 22232 41788 22524 42080 sw
tri 22524 41788 22816 42080 ne
rect 22816 41902 26664 42080
tri 26664 41902 26946 42184 sw
tri 26946 41902 27228 42184 ne
rect 27228 41929 31148 42184
tri 31148 41929 31445 42226 sw
tri 31445 41929 31742 42226 ne
rect 31742 42151 33211 42226
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42151 35480 42440
rect 31742 41929 33500 42151
rect 27228 41902 31445 41929
rect 22816 41788 26946 41902
rect 21648 41496 22524 41788
tri 22524 41496 22816 41788 sw
tri 22816 41496 23108 41788 ne
rect 23108 41620 26946 41788
tri 26946 41620 27228 41902 sw
tri 27228 41620 27510 41902 ne
rect 27510 41731 31445 41902
tri 31445 41731 31643 41929 sw
tri 31742 41731 31940 41929 ne
rect 31940 41862 33500 41929
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 42150 35480 42151
tri 35480 42150 35770 42440 sw
tri 35770 42150 36060 42440 ne
rect 36060 42438 39722 42440
tri 39722 42438 40016 42732 sw
tri 40016 42438 40310 42732 ne
rect 40310 42444 44260 42732
tri 44260 42444 44548 42732 sw
tri 44548 42444 44836 42732 ne
rect 44836 42579 48648 42732
tri 48648 42579 48945 42876 sw
tri 48945 42579 49242 42876 ne
rect 49242 42687 53085 42876
tri 53085 42687 53378 42980 sw
tri 53378 42687 53671 42980 ne
rect 53671 42800 55246 42980
tri 55246 42800 55538 43092 sw
tri 55538 42800 55830 43092 ne
rect 55830 42887 57436 43092
tri 57436 42887 57723 43174 sw
tri 57723 42887 58010 43174 ne
rect 58010 42887 70613 43174
rect 55830 42800 57723 42887
rect 53671 42687 55538 42800
rect 49242 42579 53378 42687
rect 44836 42444 48945 42579
rect 40310 42438 44548 42444
rect 36060 42150 40016 42438
rect 34078 41910 35770 42150
tri 35770 41910 36010 42150 sw
tri 36060 41910 36300 42150 ne
rect 36300 42144 40016 42150
tri 40016 42144 40310 42438 sw
tri 40310 42144 40604 42438 ne
rect 40604 42264 44548 42438
tri 44548 42264 44728 42444 sw
tri 44836 42264 45016 42444 ne
rect 45016 42282 48945 42444
tri 48945 42282 49242 42579 sw
tri 49242 42282 49539 42579 ne
rect 49539 42394 53378 42579
tri 53378 42394 53671 42687 sw
tri 53671 42394 53964 42687 ne
rect 53964 42600 55538 42687
tri 55538 42600 55738 42800 sw
tri 55830 42600 56030 42800 ne
rect 56030 42600 57723 42800
tri 57723 42600 58010 42887 sw
tri 58010 42800 58097 42887 ne
rect 58097 42875 70613 42887
rect 70669 42875 71000 45739
rect 58097 42800 71000 42875
rect 53964 42394 55738 42600
rect 49539 42282 53671 42394
rect 45016 42264 49242 42282
rect 40604 42144 44728 42264
rect 36300 41910 40310 42144
rect 34078 41862 36010 41910
rect 31940 41731 33789 41862
rect 27510 41620 31643 41731
rect 23108 41496 27228 41620
rect 21648 41204 22816 41496
tri 22816 41204 23108 41496 sw
tri 23108 41204 23400 41496 ne
rect 23400 41338 27228 41496
tri 27228 41338 27510 41620 sw
tri 27510 41338 27792 41620 ne
rect 27792 41434 31643 41620
tri 31643 41434 31940 41731 sw
tri 31940 41434 32237 41731 ne
rect 32237 41573 33789 41731
tri 33789 41573 34078 41862 sw
tri 34078 41573 34367 41862 ne
rect 34367 41620 36010 41862
tri 36010 41620 36300 41910 sw
tri 36300 41620 36590 41910 ne
rect 36590 41850 40310 41910
tri 40310 41850 40604 42144 sw
tri 40604 41850 40898 42144 ne
rect 40898 41976 44728 42144
tri 44728 41976 45016 42264 sw
tri 45016 41976 45304 42264 ne
rect 45304 41985 49242 42264
tri 49242 41985 49539 42282 sw
tri 49539 41985 49836 42282 ne
rect 49836 42101 53671 42282
tri 53671 42101 53964 42394 sw
tri 53964 42101 54257 42394 ne
rect 54257 42308 55738 42394
tri 55738 42308 56030 42600 sw
tri 56030 42308 56322 42600 ne
rect 56322 42497 71000 42600
rect 56322 42308 70613 42497
rect 54257 42101 56030 42308
rect 49836 41985 53964 42101
rect 45304 41976 49539 41985
rect 40898 41850 45016 41976
rect 36590 41620 40604 41850
rect 34367 41573 36300 41620
rect 32237 41434 34078 41573
rect 27792 41338 31940 41434
rect 23400 41204 27510 41338
rect 21648 40924 23108 41204
tri 23108 40924 23388 41204 sw
tri 23400 40924 23680 41204 ne
rect 23680 41056 27510 41204
tri 27510 41056 27792 41338 sw
tri 27792 41056 28074 41338 ne
rect 28074 41137 31940 41338
tri 31940 41137 32237 41434 sw
tri 32237 41137 32534 41434 ne
rect 32534 41297 34078 41434
tri 34078 41297 34354 41573 sw
tri 34367 41297 34643 41573 ne
rect 34643 41330 36300 41573
tri 36300 41330 36590 41620 sw
tri 36590 41330 36880 41620 ne
rect 36880 41556 40604 41620
tri 40604 41556 40898 41850 sw
tri 40898 41556 41192 41850 ne
rect 41192 41688 45016 41850
tri 45016 41688 45304 41976 sw
tri 45304 41688 45592 41976 ne
rect 45592 41688 49539 41976
tri 49539 41688 49836 41985 sw
tri 49836 41688 50133 41985 ne
rect 50133 41879 53964 41985
tri 53964 41879 54186 42101 sw
tri 54257 41879 54479 42101 ne
rect 54479 42016 56030 42101
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 70613 42308
rect 54479 41879 56322 42016
rect 50133 41688 54186 41879
rect 41192 41556 45304 41688
rect 36880 41330 40898 41556
rect 34643 41297 36590 41330
rect 32534 41137 34354 41297
rect 28074 41056 32237 41137
rect 23680 40924 27792 41056
rect 21648 40632 23388 40924
tri 23388 40632 23680 40924 sw
tri 23680 40632 23972 40924 ne
rect 23972 40774 27792 40924
tri 27792 40774 28074 41056 sw
tri 28074 40774 28356 41056 ne
rect 28356 40840 32237 41056
tri 32237 40840 32534 41137 sw
tri 32534 40840 32831 41137 ne
rect 32831 41129 34354 41137
tri 34354 41129 34522 41297 sw
tri 34643 41129 34811 41297 ne
rect 34811 41129 36590 41297
rect 32831 40840 34522 41129
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 41040 36590 41129
tri 36590 41040 36880 41330 sw
tri 36880 41040 37170 41330 ne
rect 37170 41262 40898 41330
tri 40898 41262 41192 41556 sw
tri 41192 41262 41486 41556 ne
rect 41486 41400 45304 41556
tri 45304 41400 45592 41688 sw
tri 45592 41400 45880 41688 ne
rect 45880 41400 49836 41688
rect 41486 41262 45592 41400
rect 37170 41040 41192 41262
rect 35100 40840 36880 41040
rect 28356 40774 32534 40840
rect 23972 40632 28074 40774
rect 21648 40340 23680 40632
tri 23680 40340 23972 40632 sw
tri 23972 40340 24264 40632 ne
rect 24264 40492 28074 40632
tri 28074 40492 28356 40774 sw
tri 28356 40492 28638 40774 ne
rect 28638 40543 32534 40774
tri 32534 40543 32831 40840 sw
tri 32831 40543 33128 40840 ne
rect 33128 40749 34811 40840
tri 34811 40749 34902 40840 sw
tri 35100 40749 35191 40840 ne
rect 35191 40750 36880 40840
tri 36880 40750 37170 41040 sw
tri 37170 40750 37460 41040 ne
rect 37460 41002 41192 41040
tri 41192 41002 41452 41262 sw
tri 41486 41002 41746 41262 ne
rect 41746 41112 45592 41262
tri 45592 41112 45880 41400 sw
tri 45880 41112 46168 41400 ne
rect 46168 41391 49836 41400
tri 49836 41391 50133 41688 sw
tri 50133 41391 50430 41688 ne
rect 50430 41586 54186 41688
tri 54186 41586 54479 41879 sw
tri 54479 41586 54772 41879 ne
rect 54772 41784 56322 41879
tri 56322 41784 56554 42016 sw
tri 56614 41784 56846 42016 ne
rect 56846 41784 70613 42016
rect 54772 41586 56554 41784
rect 50430 41391 54479 41586
rect 46168 41238 50133 41391
tri 50133 41238 50286 41391 sw
tri 50430 41238 50583 41391 ne
rect 50583 41293 54479 41391
tri 54479 41293 54772 41586 sw
tri 54772 41293 55065 41586 ne
rect 55065 41492 56554 41586
tri 56554 41492 56846 41784 sw
tri 56846 41492 57138 41784 ne
rect 57138 41492 70613 41784
rect 55065 41293 56846 41492
rect 50583 41238 54772 41293
rect 46168 41112 50286 41238
rect 41746 41002 45880 41112
rect 37460 40750 41452 41002
rect 35191 40749 37170 40750
rect 33128 40543 34902 40749
rect 28638 40492 32831 40543
rect 24264 40340 28356 40492
rect 21648 40048 23972 40340
tri 23972 40048 24264 40340 sw
tri 24264 40048 24556 40340 ne
rect 24556 40210 28356 40340
tri 28356 40210 28638 40492 sw
tri 28638 40210 28920 40492 ne
rect 28920 40246 32831 40492
tri 32831 40246 33128 40543 sw
tri 33128 40246 33425 40543 ne
rect 33425 40460 34902 40543
tri 34902 40460 35191 40749 sw
tri 35191 40460 35480 40749 ne
rect 35480 40460 37170 40749
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40708 41452 40750
tri 41452 40708 41746 41002 sw
tri 41746 40708 42040 41002 ne
rect 42040 40824 45880 41002
tri 45880 40824 46168 41112 sw
tri 46168 40824 46456 41112 ne
rect 46456 40941 50286 41112
tri 50286 40941 50583 41238 sw
tri 50583 40941 50880 41238 ne
rect 50880 41000 54772 41238
tri 54772 41000 55065 41293 sw
tri 55065 41000 55358 41293 ne
rect 55358 41200 56846 41293
tri 56846 41200 57138 41492 sw
tri 57138 41200 57430 41492 ne
rect 57430 41297 70613 41492
rect 70669 41297 71000 42497
rect 57430 41200 71000 41297
rect 55358 41000 57138 41200
tri 57138 41000 57338 41200 sw
rect 50880 40941 55065 41000
rect 46456 40824 50583 40941
rect 42040 40708 46168 40824
rect 37750 40460 41746 40708
rect 33425 40246 35191 40460
rect 28920 40210 33128 40246
rect 24556 40048 28638 40210
rect 21648 39756 24264 40048
tri 24264 39756 24556 40048 sw
tri 24556 39756 24848 40048 ne
rect 24848 39928 28638 40048
tri 28638 39928 28920 40210 sw
tri 28920 39928 29202 40210 ne
rect 29202 39949 33128 40210
tri 33128 39949 33425 40246 sw
tri 33425 39949 33722 40246 ne
rect 33722 40171 35191 40246
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40171 37460 40460
rect 33722 39949 35480 40171
rect 29202 39928 33425 39949
rect 24848 39830 28920 39928
tri 28920 39830 29018 39928 sw
tri 29202 39830 29300 39928 ne
rect 29300 39830 33425 39928
rect 24848 39756 29018 39830
rect 21648 39464 24556 39756
tri 24556 39464 24848 39756 sw
tri 24848 39464 25140 39756 ne
rect 25140 39548 29018 39756
tri 29018 39548 29300 39830 sw
tri 29300 39548 29582 39830 ne
rect 29582 39751 33425 39830
tri 33425 39751 33623 39949 sw
tri 33722 39751 33920 39949 ne
rect 33920 39882 35480 39949
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40170 37460 40171
tri 37460 40170 37750 40460 sw
tri 37750 40170 38040 40460 ne
rect 38040 40414 41746 40460
tri 41746 40414 42040 40708 sw
tri 42040 40414 42334 40708 ne
rect 42334 40536 46168 40708
tri 46168 40536 46456 40824 sw
tri 46456 40536 46744 40824 ne
rect 46744 40644 50583 40824
tri 50583 40644 50880 40941 sw
tri 50880 40644 51177 40941 ne
rect 51177 40707 55065 40941
tri 55065 40707 55358 41000 sw
tri 55358 40707 55651 41000 ne
rect 55651 40707 71000 41000
rect 51177 40644 55358 40707
rect 46744 40536 50880 40644
rect 42334 40414 46456 40536
rect 38040 40170 42040 40414
rect 36058 39882 37750 40170
rect 33920 39751 35769 39882
rect 29582 39548 33623 39751
rect 25140 39464 29300 39548
rect 21648 39172 24848 39464
tri 24848 39172 25140 39464 sw
tri 25140 39172 25432 39464 ne
rect 25432 39266 29300 39464
tri 29300 39266 29582 39548 sw
tri 29582 39266 29864 39548 ne
rect 29864 39454 33623 39548
tri 33623 39454 33920 39751 sw
tri 33920 39454 34217 39751 ne
rect 34217 39593 35769 39751
tri 35769 39593 36058 39882 sw
tri 36058 39593 36347 39882 ne
rect 36347 39880 37750 39882
tri 37750 39880 38040 40170 sw
tri 38040 39880 38330 40170 ne
rect 38330 40120 42040 40170
tri 42040 40120 42334 40414 sw
tri 42334 40120 42628 40414 ne
rect 42628 40248 46456 40414
tri 46456 40248 46744 40536 sw
tri 46744 40248 47032 40536 ne
rect 47032 40347 50880 40536
tri 50880 40347 51177 40644 sw
tri 51177 40347 51474 40644 ne
rect 51474 40414 55358 40644
tri 55358 40414 55651 40707 sw
tri 55651 40414 55944 40707 ne
rect 55944 40414 71000 40707
rect 51474 40347 55651 40414
rect 47032 40248 51177 40347
rect 42628 40120 46744 40248
rect 38330 39880 42334 40120
rect 36347 39822 38040 39880
tri 38040 39822 38098 39880 sw
tri 38330 39822 38388 39880 ne
rect 38388 39826 42334 39880
tri 42334 39826 42628 40120 sw
tri 42628 39826 42922 40120 ne
rect 42922 39960 46744 40120
tri 46744 39960 47032 40248 sw
tri 47032 39960 47320 40248 ne
rect 47320 40050 51177 40248
tri 51177 40050 51474 40347 sw
tri 51474 40050 51771 40347 ne
rect 51771 40186 55651 40347
tri 55651 40186 55879 40414 sw
tri 55944 40186 56172 40414 ne
rect 56172 40186 71000 40414
rect 51771 40050 55879 40186
rect 47320 39960 51474 40050
rect 42922 39928 47032 39960
tri 47032 39928 47064 39960 sw
tri 47320 39928 47352 39960 ne
rect 47352 39928 51474 39960
rect 42922 39826 47064 39928
rect 38388 39822 42628 39826
rect 36347 39593 38098 39822
rect 34217 39454 36058 39593
rect 29864 39266 33920 39454
rect 25432 39172 29582 39266
rect 21648 39004 25140 39172
tri 25140 39004 25308 39172 sw
tri 25432 39004 25600 39172 ne
rect 25600 39004 29582 39172
rect 21648 38712 25308 39004
tri 25308 38712 25600 39004 sw
tri 25600 38712 25892 39004 ne
rect 25892 38984 29582 39004
tri 29582 38984 29864 39266 sw
tri 29864 38984 30146 39266 ne
rect 30146 39157 33920 39266
tri 33920 39157 34217 39454 sw
tri 34217 39157 34514 39454 ne
rect 34514 39332 36058 39454
tri 36058 39332 36319 39593 sw
tri 36347 39332 36608 39593 ne
rect 36608 39532 38098 39593
tri 38098 39532 38388 39822 sw
tri 38388 39532 38678 39822 ne
rect 38678 39532 42628 39822
tri 42628 39532 42922 39826 sw
tri 42922 39532 43216 39826 ne
rect 43216 39640 47064 39826
tri 47064 39640 47352 39928 sw
tri 47352 39640 47640 39928 ne
rect 47640 39753 51474 39928
tri 51474 39753 51771 40050 sw
tri 51771 39753 52068 40050 ne
rect 52068 39893 55879 40050
tri 55879 39893 56172 40186 sw
tri 56172 39893 56465 40186 ne
rect 56465 39893 71000 40186
rect 52068 39753 56172 39893
rect 47640 39640 51771 39753
rect 43216 39532 47352 39640
rect 36608 39332 38388 39532
rect 34514 39157 36319 39332
rect 30146 38984 34217 39157
rect 25892 38712 29864 38984
rect 21648 38420 25600 38712
tri 25600 38420 25892 38712 sw
tri 25892 38420 26184 38712 ne
rect 26184 38702 29864 38712
tri 29864 38702 30146 38984 sw
tri 30146 38702 30428 38984 ne
rect 30428 38860 34217 38984
tri 34217 38860 34514 39157 sw
tri 34514 38860 34811 39157 ne
rect 34811 39149 36319 39157
tri 36319 39149 36502 39332 sw
tri 36608 39149 36791 39332 ne
rect 36791 39242 38388 39332
tri 38388 39242 38678 39532 sw
tri 38678 39242 38968 39532 ne
rect 38968 39242 42922 39532
rect 36791 39149 38678 39242
rect 34811 38860 36502 39149
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 39060 38678 39149
tri 38678 39060 38860 39242 sw
tri 38968 39060 39150 39242 ne
rect 39150 39238 42922 39242
tri 42922 39238 43216 39532 sw
tri 43216 39238 43510 39532 ne
rect 43510 39352 47352 39532
tri 47352 39352 47640 39640 sw
tri 47640 39352 47928 39640 ne
rect 47928 39456 51771 39640
tri 51771 39456 52068 39753 sw
tri 52068 39456 52365 39753 ne
rect 52365 39600 56172 39753
tri 56172 39600 56465 39893 sw
tri 56465 39600 56758 39893 ne
rect 56758 39600 71000 39893
rect 52365 39456 56465 39600
rect 47928 39352 52068 39456
rect 43510 39238 47640 39352
rect 39150 39076 43216 39238
tri 43216 39076 43378 39238 sw
tri 43510 39076 43672 39238 ne
rect 43672 39076 47640 39238
rect 39150 39060 43378 39076
rect 37080 38860 38860 39060
rect 30428 38702 34514 38860
rect 26184 38420 30146 38702
tri 30146 38420 30428 38702 sw
tri 30428 38420 30710 38702 ne
rect 30710 38563 34514 38702
tri 34514 38563 34811 38860 sw
tri 34811 38563 35108 38860 ne
rect 35108 38769 36791 38860
tri 36791 38769 36882 38860 sw
tri 37080 38769 37171 38860 ne
rect 37171 38770 38860 38860
tri 38860 38770 39150 39060 sw
tri 39150 38770 39440 39060 ne
rect 39440 38782 43378 39060
tri 43378 38782 43672 39076 sw
tri 43672 38782 43966 39076 ne
rect 43966 39064 47640 39076
tri 47640 39064 47928 39352 sw
tri 47928 39064 48216 39352 ne
rect 48216 39159 52068 39352
tri 52068 39159 52365 39456 sw
tri 52365 39159 52662 39456 ne
rect 52662 39400 56465 39456
tri 56465 39400 56665 39600 sw
rect 52662 39332 71000 39400
rect 52662 39159 70613 39332
rect 48216 39064 52365 39159
rect 43966 38782 47928 39064
rect 39440 38770 43672 38782
rect 37171 38769 39150 38770
rect 35108 38563 36882 38769
rect 30710 38420 34811 38563
tri 21648 34176 25892 38420 ne
tri 25892 38128 26184 38420 sw
tri 26184 38128 26476 38420 ne
rect 26476 38138 30428 38420
tri 30428 38138 30710 38420 sw
tri 30710 38138 30992 38420 ne
rect 30992 38266 34811 38420
tri 34811 38266 35108 38563 sw
tri 35108 38266 35405 38563 ne
rect 35405 38480 36882 38563
tri 36882 38480 37171 38769 sw
tri 37171 38480 37460 38769 ne
rect 37460 38480 39150 38769
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38488 43672 38770
tri 43672 38488 43966 38782 sw
tri 43966 38488 44260 38782 ne
rect 44260 38776 47928 38782
tri 47928 38776 48216 39064 sw
tri 48216 38776 48504 39064 ne
rect 48504 38929 52365 39064
tri 52365 38929 52595 39159 sw
tri 52662 38929 52892 39159 ne
rect 52892 38929 70613 39159
rect 48504 38776 52595 38929
rect 44260 38488 48216 38776
tri 48216 38488 48504 38776 sw
tri 48504 38488 48792 38776 ne
rect 48792 38632 52595 38776
tri 52595 38632 52892 38929 sw
tri 52892 38632 53189 38929 ne
rect 53189 38632 70613 38929
rect 48792 38488 52892 38632
rect 39730 38480 43966 38488
rect 35405 38266 37171 38480
rect 30992 38138 35108 38266
rect 26476 38128 30710 38138
rect 25892 37836 26184 38128
tri 26184 37836 26476 38128 sw
tri 26476 37836 26768 38128 ne
rect 26768 37940 30710 38128
tri 30710 37940 30908 38138 sw
tri 30992 37940 31190 38138 ne
rect 31190 37969 35108 38138
tri 35108 37969 35405 38266 sw
tri 35405 37969 35702 38266 ne
rect 35702 38191 37171 38266
tri 37171 38191 37460 38480 sw
tri 37460 38191 37749 38480 ne
rect 37749 38191 39440 38480
rect 35702 37969 37460 38191
rect 31190 37940 35405 37969
rect 26768 37836 30908 37940
rect 25892 37544 26476 37836
tri 26476 37544 26768 37836 sw
tri 26768 37544 27060 37836 ne
rect 27060 37658 30908 37836
tri 30908 37658 31190 37940 sw
tri 31190 37658 31472 37940 ne
rect 31472 37771 35405 37940
tri 35405 37771 35603 37969 sw
tri 35702 37771 35900 37969 ne
rect 35900 37902 37460 37969
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 38190 39440 38191
tri 39440 38190 39730 38480 sw
tri 39730 38190 40020 38480 ne
rect 40020 38194 43966 38480
tri 43966 38194 44260 38488 sw
tri 44260 38194 44554 38488 ne
rect 44554 38200 48504 38488
tri 48504 38200 48792 38488 sw
tri 48792 38200 49080 38488 ne
rect 49080 38335 52892 38488
tri 52892 38335 53189 38632 sw
tri 53189 38335 53486 38632 ne
rect 53486 38335 70613 38632
rect 49080 38200 53189 38335
rect 44554 38194 48792 38200
rect 40020 38190 44260 38194
rect 38038 37902 39730 38190
rect 35900 37771 37749 37902
rect 31472 37658 35603 37771
rect 27060 37544 31190 37658
rect 25892 37252 26768 37544
tri 26768 37252 27060 37544 sw
tri 27060 37252 27352 37544 ne
rect 27352 37376 31190 37544
tri 31190 37376 31472 37658 sw
tri 31472 37376 31754 37658 ne
rect 31754 37474 35603 37658
tri 35603 37474 35900 37771 sw
tri 35900 37474 36197 37771 ne
rect 36197 37613 37749 37771
tri 37749 37613 38038 37902 sw
tri 38038 37613 38327 37902 ne
rect 38327 37900 39730 37902
tri 39730 37900 40020 38190 sw
tri 40020 37900 40310 38190 ne
rect 40310 37900 44260 38190
tri 44260 37900 44554 38194 sw
tri 44554 37900 44848 38194 ne
rect 44848 38020 48792 38194
tri 48792 38020 48972 38200 sw
tri 49080 38020 49260 38200 ne
rect 49260 38038 53189 38200
tri 53189 38038 53486 38335 sw
tri 53486 38038 53783 38335 ne
rect 53783 38038 70613 38335
rect 49260 38020 53486 38038
rect 44848 37900 48972 38020
rect 38327 37666 40020 37900
tri 40020 37666 40254 37900 sw
tri 40310 37666 40544 37900 ne
rect 40544 37666 44554 37900
rect 38327 37613 40254 37666
rect 36197 37474 38038 37613
rect 31754 37376 35900 37474
rect 27352 37252 31472 37376
rect 25892 36960 27060 37252
tri 27060 36960 27352 37252 sw
tri 27352 36960 27644 37252 ne
rect 27644 37094 31472 37252
tri 31472 37094 31754 37376 sw
tri 31754 37094 32036 37376 ne
rect 32036 37177 35900 37376
tri 35900 37177 36197 37474 sw
tri 36197 37177 36494 37474 ne
rect 36494 37458 38038 37474
tri 38038 37458 38193 37613 sw
tri 38327 37458 38482 37613 ne
rect 38482 37458 40254 37613
rect 36494 37177 38193 37458
rect 32036 37094 36197 37177
rect 27644 36960 31754 37094
rect 25892 36680 27352 36960
tri 27352 36680 27632 36960 sw
tri 27644 36680 27924 36960 ne
rect 27924 36812 31754 36960
tri 31754 36812 32036 37094 sw
tri 32036 36812 32318 37094 ne
rect 32318 36880 36197 37094
tri 36197 36880 36494 37177 sw
tri 36494 36880 36791 37177 ne
rect 36791 37169 38193 37177
tri 38193 37169 38482 37458 sw
tri 38482 37169 38771 37458 ne
rect 38771 37376 40254 37458
tri 40254 37376 40544 37666 sw
tri 40544 37376 40834 37666 ne
rect 40834 37606 44554 37666
tri 44554 37606 44848 37900 sw
tri 44848 37606 45142 37900 ne
rect 45142 37732 48972 37900
tri 48972 37732 49260 38020 sw
tri 49260 37732 49548 38020 ne
rect 49548 37741 53486 38020
tri 53486 37741 53783 38038 sw
tri 53783 37741 54080 38038 ne
rect 54080 37741 70613 38038
rect 49548 37732 53783 37741
rect 45142 37606 49260 37732
rect 40834 37376 44848 37606
rect 38771 37169 40544 37376
rect 36791 36880 38482 37169
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 37086 40544 37169
tri 40544 37086 40834 37376 sw
tri 40834 37086 41124 37376 ne
rect 41124 37312 44848 37376
tri 44848 37312 45142 37606 sw
tri 45142 37312 45436 37606 ne
rect 45436 37444 49260 37606
tri 49260 37444 49548 37732 sw
tri 49548 37444 49836 37732 ne
rect 49836 37444 53783 37732
tri 53783 37444 54080 37741 sw
tri 54080 37444 54377 37741 ne
rect 54377 37444 70613 37741
rect 45436 37312 49548 37444
rect 41124 37086 45142 37312
rect 39060 36880 40834 37086
tri 40834 36880 41040 37086 sw
tri 41124 36880 41330 37086 ne
rect 41330 37018 45142 37086
tri 45142 37018 45436 37312 sw
tri 45436 37018 45730 37312 ne
rect 45730 37156 49548 37312
tri 49548 37156 49836 37444 sw
tri 49836 37156 50124 37444 ne
rect 50124 37156 54080 37444
rect 45730 37018 49836 37156
rect 41330 36880 45436 37018
rect 32318 36812 36494 36880
rect 27924 36680 32036 36812
rect 25892 36388 27632 36680
tri 27632 36388 27924 36680 sw
tri 27924 36388 28216 36680 ne
rect 28216 36530 32036 36680
tri 32036 36530 32318 36812 sw
tri 32318 36530 32600 36812 ne
rect 32600 36583 36494 36812
tri 36494 36583 36791 36880 sw
tri 36791 36583 37088 36880 ne
rect 37088 36789 38771 36880
tri 38771 36789 38862 36880 sw
tri 39060 36789 39151 36880 ne
rect 39151 36790 41040 36880
tri 41040 36790 41130 36880 sw
tri 41330 36790 41420 36880 ne
rect 41420 36790 45436 36880
rect 39151 36789 41130 36790
rect 37088 36583 38862 36789
rect 32600 36530 36791 36583
rect 28216 36388 32318 36530
rect 25892 36096 27924 36388
tri 27924 36096 28216 36388 sw
tri 28216 36096 28508 36388 ne
rect 28508 36248 32318 36388
tri 32318 36248 32600 36530 sw
tri 32600 36248 32882 36530 ne
rect 32882 36286 36791 36530
tri 36791 36286 37088 36583 sw
tri 37088 36286 37385 36583 ne
rect 37385 36500 38862 36583
tri 38862 36500 39151 36789 sw
tri 39151 36500 39440 36789 ne
rect 39440 36500 41130 36789
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36758 45436 36790
tri 45436 36758 45696 37018 sw
tri 45730 36758 45990 37018 ne
rect 45990 36868 49836 37018
tri 49836 36868 50124 37156 sw
tri 50124 36868 50412 37156 ne
rect 50412 37147 54080 37156
tri 54080 37147 54377 37444 sw
tri 54377 37147 54674 37444 ne
rect 54674 37147 70613 37444
rect 50412 36994 54377 37147
tri 54377 36994 54530 37147 sw
tri 54674 36994 54827 37147 ne
rect 54827 36994 70613 37147
rect 50412 36868 54530 36994
rect 45990 36758 50124 36868
rect 41710 36500 45696 36758
rect 37385 36286 39151 36500
rect 32882 36248 37088 36286
rect 28508 36096 32600 36248
rect 25892 35804 28216 36096
tri 28216 35804 28508 36096 sw
tri 28508 35804 28800 36096 ne
rect 28800 35966 32600 36096
tri 32600 35966 32882 36248 sw
tri 32882 35966 33164 36248 ne
rect 33164 35989 37088 36248
tri 37088 35989 37385 36286 sw
tri 37385 35989 37682 36286 ne
rect 37682 36211 39151 36286
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36211 41420 36500
rect 37682 35989 39440 36211
rect 33164 35966 37385 35989
rect 28800 35804 32882 35966
rect 25892 35512 28508 35804
tri 28508 35512 28800 35804 sw
tri 28800 35512 29092 35804 ne
rect 29092 35684 32882 35804
tri 32882 35684 33164 35966 sw
tri 33164 35684 33446 35966 ne
rect 33446 35791 37385 35966
tri 37385 35791 37583 35989 sw
tri 37682 35791 37880 35989 ne
rect 37880 35922 39440 35989
tri 39440 35922 39729 36211 sw
tri 39729 35922 40018 36211 ne
rect 40018 36210 41420 36211
tri 41420 36210 41710 36500 sw
tri 41710 36210 42000 36500 ne
rect 42000 36464 45696 36500
tri 45696 36464 45990 36758 sw
tri 45990 36464 46284 36758 ne
rect 46284 36580 50124 36758
tri 50124 36580 50412 36868 sw
tri 50412 36580 50700 36868 ne
rect 50700 36697 54530 36868
tri 54530 36697 54827 36994 sw
tri 54827 36697 55124 36994 ne
rect 55124 36697 70613 36994
rect 50700 36580 54827 36697
rect 46284 36464 50412 36580
rect 42000 36210 45990 36464
rect 40018 35922 41710 36210
rect 37880 35791 39729 35922
rect 33446 35684 37583 35791
rect 29092 35586 33164 35684
tri 33164 35586 33262 35684 sw
tri 33446 35586 33544 35684 ne
rect 33544 35586 37583 35684
rect 29092 35512 33262 35586
rect 25892 35220 28800 35512
tri 28800 35220 29092 35512 sw
tri 29092 35220 29384 35512 ne
rect 29384 35304 33262 35512
tri 33262 35304 33544 35586 sw
tri 33544 35304 33826 35586 ne
rect 33826 35494 37583 35586
tri 37583 35494 37880 35791 sw
tri 37880 35494 38177 35791 ne
rect 38177 35633 39729 35791
tri 39729 35633 40018 35922 sw
tri 40018 35633 40307 35922 ne
rect 40307 35920 41710 35922
tri 41710 35920 42000 36210 sw
tri 42000 35920 42290 36210 ne
rect 42290 36170 45990 36210
tri 45990 36170 46284 36464 sw
tri 46284 36170 46578 36464 ne
rect 46578 36292 50412 36464
tri 50412 36292 50700 36580 sw
tri 50700 36292 50988 36580 ne
rect 50988 36400 54827 36580
tri 54827 36400 55124 36697 sw
tri 55124 36400 55421 36697 ne
rect 55421 36468 70613 36697
rect 70669 36468 71000 39332
rect 55421 36400 71000 36468
rect 50988 36292 55124 36400
rect 46578 36170 50700 36292
rect 42290 35920 46284 36170
rect 40307 35868 42000 35920
tri 42000 35868 42052 35920 sw
tri 42290 35868 42342 35920 ne
rect 42342 35876 46284 35920
tri 46284 35876 46578 36170 sw
tri 46578 35876 46872 36170 ne
rect 46872 36004 50700 36170
tri 50700 36004 50988 36292 sw
tri 50988 36004 51276 36292 ne
rect 51276 36200 55124 36292
tri 55124 36200 55324 36400 sw
rect 51276 36132 71000 36200
rect 51276 36004 70613 36132
rect 46872 35876 50988 36004
rect 42342 35868 46578 35876
rect 40307 35633 42052 35868
rect 38177 35494 40018 35633
rect 33826 35304 37880 35494
rect 29384 35220 33544 35304
rect 25892 34928 29092 35220
tri 29092 34928 29384 35220 sw
tri 29384 34928 29676 35220 ne
rect 29676 35022 33544 35220
tri 33544 35022 33826 35304 sw
tri 33826 35022 34108 35304 ne
rect 34108 35197 37880 35304
tri 37880 35197 38177 35494 sw
tri 38177 35197 38474 35494 ne
rect 38474 35478 40018 35494
tri 40018 35478 40173 35633 sw
tri 40307 35478 40462 35633 ne
rect 40462 35578 42052 35633
tri 42052 35578 42342 35868 sw
tri 42342 35578 42632 35868 ne
rect 42632 35582 46578 35868
tri 46578 35582 46872 35876 sw
tri 46872 35582 47166 35876 ne
rect 47166 35716 50988 35876
tri 50988 35716 51276 36004 sw
tri 51276 35716 51564 36004 ne
rect 51564 35716 70613 36004
rect 47166 35684 51276 35716
tri 51276 35684 51308 35716 sw
tri 51564 35684 51596 35716 ne
rect 51596 35684 70613 35716
rect 47166 35582 51308 35684
rect 42632 35578 46872 35582
rect 40462 35478 42342 35578
rect 38474 35197 40173 35478
rect 34108 35022 38177 35197
rect 29676 34928 33826 35022
rect 25892 34760 29384 34928
tri 29384 34760 29552 34928 sw
tri 29676 34760 29844 34928 ne
rect 29844 34760 33826 34928
rect 25892 34468 29552 34760
tri 29552 34468 29844 34760 sw
tri 29844 34468 30136 34760 ne
rect 30136 34740 33826 34760
tri 33826 34740 34108 35022 sw
tri 34108 34740 34390 35022 ne
rect 34390 34900 38177 35022
tri 38177 34900 38474 35197 sw
tri 38474 34900 38771 35197 ne
rect 38771 35189 40173 35197
tri 40173 35189 40462 35478 sw
tri 40462 35189 40751 35478 ne
rect 40751 35288 42342 35478
tri 42342 35288 42632 35578 sw
tri 42632 35288 42922 35578 ne
rect 42922 35288 46872 35578
tri 46872 35288 47166 35582 sw
tri 47166 35288 47460 35582 ne
rect 47460 35396 51308 35582
tri 51308 35396 51596 35684 sw
tri 51596 35396 51884 35684 ne
rect 51884 35396 70613 35684
rect 47460 35288 51596 35396
rect 40751 35189 42632 35288
rect 38771 34900 40462 35189
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42632 35189
tri 42632 34998 42922 35288 sw
tri 42922 34998 43212 35288 ne
rect 43212 34998 47166 35288
rect 41040 34900 42922 34998
rect 34390 34740 38474 34900
rect 30136 34468 34108 34740
rect 25892 34176 29844 34468
tri 29844 34176 30136 34468 sw
tri 30136 34176 30428 34468 ne
rect 30428 34458 34108 34468
tri 34108 34458 34390 34740 sw
tri 34390 34458 34672 34740 ne
rect 34672 34603 38474 34740
tri 38474 34603 38771 34900 sw
tri 38771 34603 39068 34900 ne
rect 39068 34809 40751 34900
tri 40751 34809 40842 34900 sw
tri 41040 34809 41131 34900 ne
rect 41131 34810 42922 34900
tri 42922 34810 43110 34998 sw
tri 43212 34810 43400 34998 ne
rect 43400 34994 47166 34998
tri 47166 34994 47460 35288 sw
tri 47460 34994 47754 35288 ne
rect 47754 35108 51596 35288
tri 51596 35108 51884 35396 sw
tri 51884 35108 52172 35396 ne
rect 52172 35108 70613 35396
rect 47754 34994 51884 35108
rect 43400 34832 47460 34994
tri 47460 34832 47622 34994 sw
tri 47754 34832 47916 34994 ne
rect 47916 34832 51884 34994
rect 43400 34810 47622 34832
rect 41131 34809 43110 34810
rect 39068 34603 40842 34809
rect 34672 34458 38771 34603
rect 30428 34176 34390 34458
tri 34390 34176 34672 34458 sw
tri 34672 34176 34954 34458 ne
rect 34954 34306 38771 34458
tri 38771 34306 39068 34603 sw
tri 39068 34306 39365 34603 ne
rect 39365 34520 40842 34603
tri 40842 34520 41131 34809 sw
tri 41131 34520 41420 34809 ne
rect 41420 34520 43110 34809
tri 43110 34520 43400 34810 sw
tri 43400 34520 43690 34810 ne
rect 43690 34538 47622 34810
tri 47622 34538 47916 34832 sw
tri 47916 34538 48210 34832 ne
rect 48210 34820 51884 34832
tri 51884 34820 52172 35108 sw
tri 52172 34820 52460 35108 ne
rect 52460 34820 70613 35108
rect 48210 34538 52172 34820
rect 43690 34520 47916 34538
rect 39365 34306 41131 34520
rect 34954 34176 39068 34306
tri 25892 29932 30136 34176 ne
tri 30136 33884 30428 34176 sw
tri 30428 33884 30720 34176 ne
rect 30720 33894 34672 34176
tri 34672 33894 34954 34176 sw
tri 34954 33894 35236 34176 ne
rect 35236 34009 39068 34176
tri 39068 34009 39365 34306 sw
tri 39365 34009 39662 34306 ne
rect 39662 34231 41131 34306
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34244 43400 34520
tri 43400 34244 43676 34520 sw
tri 43690 34244 43966 34520 ne
rect 43966 34244 47916 34520
tri 47916 34244 48210 34538 sw
tri 48210 34244 48504 34538 ne
rect 48504 34532 52172 34538
tri 52172 34532 52460 34820 sw
tri 52460 34532 52748 34820 ne
rect 52748 34532 70613 34820
rect 48504 34244 52460 34532
tri 52460 34244 52748 34532 sw
tri 52748 34244 53036 34532 ne
rect 53036 34244 70613 34532
rect 41709 34231 43676 34244
rect 39662 34009 41420 34231
rect 35236 33894 39365 34009
rect 30720 33884 34954 33894
rect 30136 33592 30428 33884
tri 30428 33592 30720 33884 sw
tri 30720 33592 31012 33884 ne
rect 31012 33696 34954 33884
tri 34954 33696 35152 33894 sw
tri 35236 33696 35434 33894 ne
rect 35434 33811 39365 33894
tri 39365 33811 39563 34009 sw
tri 39662 33811 39860 34009 ne
rect 39860 33942 41420 34009
tri 41420 33942 41709 34231 sw
tri 41709 33942 41998 34231 ne
rect 41998 33954 43676 34231
tri 43676 33954 43966 34244 sw
tri 43966 33954 44256 34244 ne
rect 44256 33954 48210 34244
rect 41998 33942 43966 33954
rect 39860 33811 41709 33942
rect 35434 33696 39563 33811
rect 31012 33592 35152 33696
rect 30136 33300 30720 33592
tri 30720 33300 31012 33592 sw
tri 31012 33300 31304 33592 ne
rect 31304 33414 35152 33592
tri 35152 33414 35434 33696 sw
tri 35434 33414 35716 33696 ne
rect 35716 33514 39563 33696
tri 39563 33514 39860 33811 sw
tri 39860 33514 40157 33811 ne
rect 40157 33653 41709 33811
tri 41709 33653 41998 33942 sw
tri 41998 33653 42287 33942 ne
rect 42287 33664 43966 33942
tri 43966 33664 44256 33954 sw
tri 44256 33664 44546 33954 ne
rect 44546 33950 48210 33954
tri 48210 33950 48504 34244 sw
tri 48504 33950 48798 34244 ne
rect 48798 33956 52748 34244
tri 52748 33956 53036 34244 sw
tri 53036 33956 53324 34244 ne
rect 53324 33956 70613 34244
rect 48798 33950 53036 33956
rect 44546 33664 48504 33950
rect 42287 33653 44256 33664
rect 40157 33514 41998 33653
rect 35716 33414 39860 33514
rect 31304 33300 35434 33414
rect 30136 33008 31012 33300
tri 31012 33008 31304 33300 sw
tri 31304 33008 31596 33300 ne
rect 31596 33132 35434 33300
tri 35434 33132 35716 33414 sw
tri 35716 33132 35998 33414 ne
rect 35998 33217 39860 33414
tri 39860 33217 40157 33514 sw
tri 40157 33217 40454 33514 ne
rect 40454 33498 41998 33514
tri 41998 33498 42153 33653 sw
tri 42287 33498 42442 33653 ne
rect 42442 33498 44256 33653
rect 40454 33217 42153 33498
rect 35998 33132 40157 33217
rect 31596 33008 35716 33132
rect 30136 32716 31304 33008
tri 31304 32716 31596 33008 sw
tri 31596 32716 31888 33008 ne
rect 31888 32850 35716 33008
tri 35716 32850 35998 33132 sw
tri 35998 32850 36280 33132 ne
rect 36280 32920 40157 33132
tri 40157 32920 40454 33217 sw
tri 40454 32920 40751 33217 ne
rect 40751 33209 42153 33217
tri 42153 33209 42442 33498 sw
tri 42442 33209 42731 33498 ne
rect 42731 33422 44256 33498
tri 44256 33422 44498 33664 sw
tri 44546 33422 44788 33664 ne
rect 44788 33656 48504 33664
tri 48504 33656 48798 33950 sw
tri 48798 33656 49092 33950 ne
rect 49092 33776 53036 33950
tri 53036 33776 53216 33956 sw
tri 53324 33776 53504 33956 ne
rect 53504 33776 70613 33956
rect 49092 33656 53216 33776
rect 44788 33422 48798 33656
rect 42731 33209 44498 33422
rect 40751 32920 42442 33209
tri 42442 32920 42731 33209 sw
tri 42731 32920 43020 33209 ne
rect 43020 33132 44498 33209
tri 44498 33132 44788 33422 sw
tri 44788 33132 45078 33422 ne
rect 45078 33362 48798 33422
tri 48798 33362 49092 33656 sw
tri 49092 33362 49386 33656 ne
rect 49386 33488 53216 33656
tri 53216 33488 53504 33776 sw
tri 53504 33488 53792 33776 ne
rect 53792 33488 70613 33776
rect 49386 33362 53504 33488
rect 45078 33132 49092 33362
rect 43020 32920 44788 33132
rect 36280 32850 40454 32920
rect 31888 32716 35998 32850
rect 30136 32436 31596 32716
tri 31596 32436 31876 32716 sw
tri 31888 32436 32168 32716 ne
rect 32168 32568 35998 32716
tri 35998 32568 36280 32850 sw
tri 36280 32568 36562 32850 ne
rect 36562 32623 40454 32850
tri 40454 32623 40751 32920 sw
tri 40751 32623 41048 32920 ne
rect 41048 32829 42731 32920
tri 42731 32829 42822 32920 sw
tri 43020 32829 43111 32920 ne
rect 43111 32842 44788 32920
tri 44788 32842 45078 33132 sw
tri 45078 32842 45368 33132 ne
rect 45368 33068 49092 33132
tri 49092 33068 49386 33362 sw
tri 49386 33068 49680 33362 ne
rect 49680 33200 53504 33362
tri 53504 33200 53792 33488 sw
tri 53792 33200 54080 33488 ne
rect 54080 33268 70613 33488
rect 70669 33268 71000 36132
rect 54080 33200 71000 33268
rect 49680 33068 53792 33200
rect 45368 32842 49386 33068
rect 43111 32830 45078 32842
tri 45078 32830 45090 32842 sw
tri 45368 32830 45380 32842 ne
rect 45380 32830 49386 32842
rect 43111 32829 45090 32830
rect 41048 32623 42822 32829
rect 36562 32568 40751 32623
rect 32168 32436 36280 32568
rect 30136 32144 31876 32436
tri 31876 32144 32168 32436 sw
tri 32168 32144 32460 32436 ne
rect 32460 32286 36280 32436
tri 36280 32286 36562 32568 sw
tri 36562 32286 36844 32568 ne
rect 36844 32326 40751 32568
tri 40751 32326 41048 32623 sw
tri 41048 32326 41345 32623 ne
rect 41345 32540 42822 32623
tri 42822 32540 43111 32829 sw
tri 43111 32540 43400 32829 ne
rect 43400 32540 45090 32829
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32774 49386 32830
tri 49386 32774 49680 33068 sw
tri 49680 32774 49974 33068 ne
rect 49974 33000 53792 33068
tri 53792 33000 53992 33200 sw
rect 49974 32920 71000 33000
rect 49974 32774 70613 32920
rect 45670 32540 49680 32774
rect 41345 32326 43111 32540
rect 36844 32286 41048 32326
rect 32460 32144 36562 32286
rect 30136 31852 32168 32144
tri 32168 31852 32460 32144 sw
tri 32460 31852 32752 32144 ne
rect 32752 32004 36562 32144
tri 36562 32004 36844 32286 sw
tri 36844 32004 37126 32286 ne
rect 37126 32029 41048 32286
tri 41048 32029 41345 32326 sw
tri 41345 32029 41642 32326 ne
rect 41642 32251 43111 32326
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32251 45380 32540
rect 41642 32029 43400 32251
rect 37126 32004 41345 32029
rect 32752 31852 36844 32004
rect 30136 31560 32460 31852
tri 32460 31560 32752 31852 sw
tri 32752 31560 33044 31852 ne
rect 33044 31722 36844 31852
tri 36844 31722 37126 32004 sw
tri 37126 31722 37408 32004 ne
rect 37408 31831 41345 32004
tri 41345 31831 41543 32029 sw
tri 41642 31831 41840 32029 ne
rect 41840 31962 43400 32029
tri 43400 31962 43689 32251 sw
tri 43689 31962 43978 32251 ne
rect 43978 32250 45380 32251
tri 45380 32250 45670 32540 sw
tri 45670 32250 45960 32540 ne
rect 45960 32514 49680 32540
tri 49680 32514 49940 32774 sw
tri 49974 32514 50234 32774 ne
rect 50234 32514 70613 32774
rect 45960 32250 49940 32514
rect 43978 31962 45670 32250
rect 41840 31831 43689 31962
rect 37408 31722 41543 31831
rect 33044 31560 37126 31722
rect 30136 31268 32752 31560
tri 32752 31268 33044 31560 sw
tri 33044 31268 33336 31560 ne
rect 33336 31440 37126 31560
tri 37126 31440 37408 31722 sw
tri 37408 31440 37690 31722 ne
rect 37690 31534 41543 31722
tri 41543 31534 41840 31831 sw
tri 41840 31534 42137 31831 ne
rect 42137 31673 43689 31831
tri 43689 31673 43978 31962 sw
tri 43978 31673 44267 31962 ne
rect 44267 31960 45670 31962
tri 45670 31960 45960 32250 sw
tri 45960 31960 46250 32250 ne
rect 46250 32220 49940 32250
tri 49940 32220 50234 32514 sw
tri 50234 32220 50528 32514 ne
rect 50528 32220 70613 32514
rect 46250 31960 50234 32220
rect 44267 31673 45960 31960
rect 42137 31534 43978 31673
rect 37690 31440 41840 31534
rect 33336 31342 37408 31440
tri 37408 31342 37506 31440 sw
tri 37690 31342 37788 31440 ne
rect 37788 31342 41840 31440
rect 33336 31268 37506 31342
rect 30136 30976 33044 31268
tri 33044 30976 33336 31268 sw
tri 33336 30976 33628 31268 ne
rect 33628 31060 37506 31268
tri 37506 31060 37788 31342 sw
tri 37788 31060 38070 31342 ne
rect 38070 31237 41840 31342
tri 41840 31237 42137 31534 sw
tri 42137 31237 42434 31534 ne
rect 42434 31518 43978 31534
tri 43978 31518 44133 31673 sw
tri 44267 31518 44422 31673 ne
rect 44422 31670 45960 31673
tri 45960 31670 46250 31960 sw
tri 46250 31670 46540 31960 ne
rect 46540 31926 50234 31960
tri 50234 31926 50528 32220 sw
tri 50528 31926 50822 32220 ne
rect 50822 31926 70613 32220
rect 46540 31670 50528 31926
rect 44422 31624 46250 31670
tri 46250 31624 46296 31670 sw
tri 46540 31624 46586 31670 ne
rect 46586 31632 50528 31670
tri 50528 31632 50822 31926 sw
tri 50822 31632 51116 31926 ne
rect 51116 31632 70613 31926
rect 46586 31624 50822 31632
rect 44422 31518 46296 31624
rect 42434 31237 44133 31518
rect 38070 31060 42137 31237
rect 33628 30976 37788 31060
rect 30136 30684 33336 30976
tri 33336 30684 33628 30976 sw
tri 33628 30684 33920 30976 ne
rect 33920 30778 37788 30976
tri 37788 30778 38070 31060 sw
tri 38070 30778 38352 31060 ne
rect 38352 30940 42137 31060
tri 42137 30940 42434 31237 sw
tri 42434 30940 42731 31237 ne
rect 42731 31229 44133 31237
tri 44133 31229 44422 31518 sw
tri 44422 31229 44711 31518 ne
rect 44711 31334 46296 31518
tri 46296 31334 46586 31624 sw
tri 46586 31334 46876 31624 ne
rect 46876 31338 50822 31624
tri 50822 31338 51116 31632 sw
tri 51116 31338 51410 31632 ne
rect 51410 31338 70613 31632
rect 46876 31334 51116 31338
rect 44711 31229 46586 31334
rect 42731 30940 44422 31229
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31044 46586 31229
tri 46586 31044 46876 31334 sw
tri 46876 31044 47166 31334 ne
rect 47166 31044 51116 31334
tri 51116 31044 51410 31338 sw
tri 51410 31044 51704 31338 ne
rect 51704 31044 70613 31338
rect 45000 30940 46876 31044
rect 38352 30778 42434 30940
rect 33920 30684 38070 30778
rect 30136 30516 33628 30684
tri 33628 30516 33796 30684 sw
tri 33920 30516 34088 30684 ne
rect 34088 30516 38070 30684
rect 30136 30224 33796 30516
tri 33796 30224 34088 30516 sw
tri 34088 30224 34380 30516 ne
rect 34380 30496 38070 30516
tri 38070 30496 38352 30778 sw
tri 38352 30496 38634 30778 ne
rect 38634 30643 42434 30778
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30849 44711 30940
tri 44711 30849 44802 30940 sw
tri 45000 30849 45091 30940 ne
rect 45091 30850 46876 30940
tri 46876 30850 47070 31044 sw
tri 47166 30850 47360 31044 ne
rect 47360 30850 51410 31044
rect 45091 30849 47070 30850
rect 43028 30643 44802 30849
rect 38634 30496 42731 30643
rect 34380 30224 38352 30496
rect 30136 29932 34088 30224
tri 34088 29932 34380 30224 sw
tri 34380 29932 34672 30224 ne
rect 34672 30214 38352 30224
tri 38352 30214 38634 30496 sw
tri 38634 30214 38916 30496 ne
rect 38916 30346 42731 30496
tri 42731 30346 43028 30643 sw
tri 43028 30346 43325 30643 ne
rect 43325 30560 44802 30643
tri 44802 30560 45091 30849 sw
tri 45091 30560 45380 30849 ne
rect 45380 30560 47070 30849
tri 47070 30560 47360 30850 sw
tri 47360 30560 47650 30850 ne
rect 47650 30750 51410 30850
tri 51410 30750 51704 31044 sw
tri 51704 30750 51998 31044 ne
rect 51998 30750 70613 31044
rect 47650 30588 51704 30750
tri 51704 30588 51866 30750 sw
tri 51998 30588 52160 30750 ne
rect 52160 30588 70613 30750
rect 47650 30560 51866 30588
rect 43325 30346 45091 30560
rect 38916 30214 43028 30346
rect 34672 29932 38634 30214
tri 38634 29932 38916 30214 sw
tri 38916 29932 39198 30214 ne
rect 39198 30049 43028 30214
tri 43028 30049 43325 30346 sw
tri 43325 30049 43622 30346 ne
rect 43622 30271 45091 30346
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30271 47360 30560
rect 43622 30049 45380 30271
rect 39198 29932 43325 30049
tri 30136 25688 34380 29932 ne
tri 34380 29640 34672 29932 sw
tri 34672 29640 34964 29932 ne
rect 34964 29650 38916 29932
tri 38916 29650 39198 29932 sw
tri 39198 29650 39480 29932 ne
rect 39480 29752 43325 29932
tri 43325 29752 43622 30049 sw
tri 43622 29752 43919 30049 ne
rect 43919 29982 45380 30049
tri 45380 29982 45669 30271 sw
tri 45669 29982 45958 30271 ne
rect 45958 30270 47360 30271
tri 47360 30270 47650 30560 sw
tri 47650 30270 47940 30560 ne
rect 47940 30294 51866 30560
tri 51866 30294 52160 30588 sw
tri 52160 30294 52454 30588 ne
rect 52454 30294 70613 30588
rect 47940 30270 52160 30294
rect 45958 30000 47650 30270
tri 47650 30000 47920 30270 sw
tri 47940 30000 48210 30270 ne
rect 48210 30000 52160 30270
tri 52160 30000 52454 30294 sw
tri 52454 30000 52748 30294 ne
rect 52748 30056 70613 30294
rect 70669 30056 71000 32920
rect 52748 30000 71000 30056
rect 45958 29982 47920 30000
rect 43919 29752 45669 29982
rect 39480 29650 43622 29752
rect 34964 29640 39198 29650
rect 34380 29348 34672 29640
tri 34672 29348 34964 29640 sw
tri 34964 29348 35256 29640 ne
rect 35256 29452 39198 29640
tri 39198 29452 39396 29650 sw
tri 39480 29452 39678 29650 ne
rect 39678 29554 43622 29650
tri 43622 29554 43820 29752 sw
tri 43919 29554 44117 29752 ne
rect 44117 29693 45669 29752
tri 45669 29693 45958 29982 sw
tri 45958 29693 46247 29982 ne
rect 46247 29710 47920 29982
tri 47920 29710 48210 30000 sw
tri 48210 29710 48500 30000 ne
rect 48500 29800 52454 30000
tri 52454 29800 52654 30000 sw
rect 48500 29752 71000 29800
rect 48500 29710 70613 29752
rect 46247 29693 48210 29710
rect 44117 29554 45958 29693
rect 39678 29452 43820 29554
rect 35256 29348 39396 29452
rect 34380 29056 34964 29348
tri 34964 29056 35256 29348 sw
tri 35256 29056 35548 29348 ne
rect 35548 29170 39396 29348
tri 39396 29170 39678 29452 sw
tri 39678 29170 39960 29452 ne
rect 39960 29257 43820 29452
tri 43820 29257 44117 29554 sw
tri 44117 29257 44414 29554 ne
rect 44414 29466 45958 29554
tri 45958 29466 46185 29693 sw
tri 46247 29466 46474 29693 ne
rect 46474 29466 48210 29693
rect 44414 29257 46185 29466
rect 39960 29170 44117 29257
rect 35548 29056 39678 29170
rect 34380 28764 35256 29056
tri 35256 28764 35548 29056 sw
tri 35548 28764 35840 29056 ne
rect 35840 28888 39678 29056
tri 39678 28888 39960 29170 sw
tri 39960 28888 40242 29170 ne
rect 40242 28960 44117 29170
tri 44117 28960 44414 29257 sw
tri 44414 28960 44711 29257 ne
rect 44711 29177 46185 29257
tri 46185 29177 46474 29466 sw
tri 46474 29177 46763 29466 ne
rect 46763 29420 48210 29466
tri 48210 29420 48500 29710 sw
tri 48500 29420 48790 29710 ne
rect 48790 29420 70613 29710
rect 46763 29178 48500 29420
tri 48500 29178 48742 29420 sw
tri 48790 29178 49032 29420 ne
rect 49032 29178 70613 29420
rect 46763 29177 48742 29178
rect 44711 28960 46474 29177
rect 40242 28888 44414 28960
rect 35840 28764 39960 28888
rect 34380 28472 35548 28764
tri 35548 28472 35840 28764 sw
tri 35840 28472 36132 28764 ne
rect 36132 28606 39960 28764
tri 39960 28606 40242 28888 sw
tri 40242 28606 40524 28888 ne
rect 40524 28663 44414 28888
tri 44414 28663 44711 28960 sw
tri 44711 28663 45008 28960 ne
rect 45008 28888 46474 28960
tri 46474 28888 46763 29177 sw
tri 46763 28888 47052 29177 ne
rect 47052 28888 48742 29177
tri 48742 28888 49032 29178 sw
tri 49032 28888 49322 29178 ne
rect 49322 28888 70613 29178
rect 45008 28869 46763 28888
tri 46763 28869 46782 28888 sw
tri 47052 28869 47071 28888 ne
rect 47071 28870 49032 28888
tri 49032 28870 49050 28888 sw
tri 49322 28870 49340 28888 ne
rect 49340 28870 70613 28888
rect 47071 28869 49050 28870
rect 45008 28663 46782 28869
rect 40524 28606 44711 28663
rect 36132 28472 40242 28606
rect 34380 28192 35840 28472
tri 35840 28192 36120 28472 sw
tri 36132 28192 36412 28472 ne
rect 36412 28324 40242 28472
tri 40242 28324 40524 28606 sw
tri 40524 28324 40806 28606 ne
rect 40806 28366 44711 28606
tri 44711 28366 45008 28663 sw
tri 45008 28366 45305 28663 ne
rect 45305 28580 46782 28663
tri 46782 28580 47071 28869 sw
tri 47071 28580 47360 28869 ne
rect 47360 28580 49050 28869
tri 49050 28580 49340 28870 sw
tri 49340 28580 49630 28870 ne
rect 49630 28580 70613 28870
rect 45305 28366 47071 28580
rect 40806 28324 45008 28366
rect 36412 28192 40524 28324
rect 34380 27900 36120 28192
tri 36120 27900 36412 28192 sw
tri 36412 27900 36704 28192 ne
rect 36704 28042 40524 28192
tri 40524 28042 40806 28324 sw
tri 40806 28042 41088 28324 ne
rect 41088 28069 45008 28324
tri 45008 28069 45305 28366 sw
tri 45305 28069 45602 28366 ne
rect 45602 28291 47071 28366
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28291 49340 28580
rect 45602 28069 47360 28291
rect 41088 28042 45305 28069
rect 36704 27900 40806 28042
rect 34380 27608 36412 27900
tri 36412 27608 36704 27900 sw
tri 36704 27608 36996 27900 ne
rect 36996 27760 40806 27900
tri 40806 27760 41088 28042 sw
tri 41088 27760 41370 28042 ne
rect 41370 27871 45305 28042
tri 45305 27871 45503 28069 sw
tri 45602 27871 45800 28069 ne
rect 45800 28002 47360 28069
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28290 49340 28291
tri 49340 28290 49630 28580 sw
tri 49630 28290 49920 28580 ne
rect 49920 28290 70613 28580
rect 47938 28002 49630 28290
rect 45800 27871 47649 28002
rect 41370 27760 45503 27871
rect 36996 27608 41088 27760
rect 34380 27316 36704 27608
tri 36704 27316 36996 27608 sw
tri 36996 27316 37288 27608 ne
rect 37288 27478 41088 27608
tri 41088 27478 41370 27760 sw
tri 41370 27478 41652 27760 ne
rect 41652 27574 45503 27760
tri 45503 27574 45800 27871 sw
tri 45800 27574 46097 27871 ne
rect 46097 27713 47649 27871
tri 47649 27713 47938 28002 sw
tri 47938 27713 48227 28002 ne
rect 48227 28000 49630 28002
tri 49630 28000 49920 28290 sw
tri 49920 28000 50210 28290 ne
rect 50210 28000 70613 28290
rect 48227 27713 49920 28000
rect 46097 27667 47938 27713
tri 47938 27667 47984 27713 sw
tri 48227 27667 48273 27713 ne
rect 48273 27710 49920 27713
tri 49920 27710 50210 28000 sw
tri 50210 27710 50500 28000 ne
rect 50500 27710 70613 28000
rect 48273 27667 50210 27710
rect 46097 27574 47984 27667
rect 41652 27478 45800 27574
rect 37288 27316 41370 27478
rect 34380 27024 36996 27316
tri 36996 27024 37288 27316 sw
tri 37288 27024 37580 27316 ne
rect 37580 27196 41370 27316
tri 41370 27196 41652 27478 sw
tri 41652 27196 41934 27478 ne
rect 41934 27277 45800 27478
tri 45800 27277 46097 27574 sw
tri 46097 27277 46394 27574 ne
rect 46394 27378 47984 27574
tri 47984 27378 48273 27667 sw
tri 48273 27378 48562 27667 ne
rect 48562 27470 50210 27667
tri 50210 27470 50450 27710 sw
tri 50500 27470 50740 27710 ne
rect 50740 27470 70613 27710
rect 48562 27378 50450 27470
rect 46394 27277 48273 27378
rect 41934 27196 46097 27277
rect 37580 27098 41652 27196
tri 41652 27098 41750 27196 sw
tri 41934 27098 42032 27196 ne
rect 42032 27098 46097 27196
rect 37580 27024 41750 27098
rect 34380 26732 37288 27024
tri 37288 26732 37580 27024 sw
tri 37580 26732 37872 27024 ne
rect 37872 26816 41750 27024
tri 41750 26816 42032 27098 sw
tri 42032 26816 42314 27098 ne
rect 42314 26980 46097 27098
tri 46097 26980 46394 27277 sw
tri 46394 26980 46691 27277 ne
rect 46691 27089 48273 27277
tri 48273 27089 48562 27378 sw
tri 48562 27089 48851 27378 ne
rect 48851 27180 50450 27378
tri 50450 27180 50740 27470 sw
tri 50740 27180 51030 27470 ne
rect 51030 27180 70613 27470
rect 48851 27089 50740 27180
rect 46691 26980 48562 27089
rect 42314 26816 46394 26980
rect 37872 26732 42032 26816
rect 34380 26440 37580 26732
tri 37580 26440 37872 26732 sw
tri 37872 26440 38164 26732 ne
rect 38164 26534 42032 26732
tri 42032 26534 42314 26816 sw
tri 42314 26534 42596 26816 ne
rect 42596 26683 46394 26816
tri 46394 26683 46691 26980 sw
tri 46691 26683 46988 26980 ne
rect 46988 26800 48562 26980
tri 48562 26800 48851 27089 sw
tri 48851 26800 49140 27089 ne
rect 49140 26890 50740 27089
tri 50740 26890 51030 27180 sw
tri 51030 26890 51320 27180 ne
rect 51320 26890 70613 27180
rect 49140 26800 51030 26890
rect 46988 26683 48851 26800
rect 42596 26534 46691 26683
rect 38164 26440 42314 26534
rect 34380 26272 37872 26440
tri 37872 26272 38040 26440 sw
tri 38164 26272 38332 26440 ne
rect 38332 26272 42314 26440
rect 34380 25980 38040 26272
tri 38040 25980 38332 26272 sw
tri 38332 25980 38624 26272 ne
rect 38624 26252 42314 26272
tri 42314 26252 42596 26534 sw
tri 42596 26252 42878 26534 ne
rect 42878 26386 46691 26534
tri 46691 26386 46988 26683 sw
tri 46988 26386 47285 26683 ne
rect 47285 26600 48851 26683
tri 48851 26600 49051 26800 sw
tri 49140 26600 49340 26800 ne
rect 49340 26600 51030 26800
tri 51030 26600 51320 26890 sw
tri 51320 26800 51410 26890 ne
rect 51410 26888 70613 26890
rect 70669 26888 71000 29752
rect 51410 26800 71000 26888
rect 47285 26386 49051 26600
rect 42878 26252 46988 26386
rect 38624 25980 42596 26252
rect 34380 25688 38332 25980
tri 38332 25688 38624 25980 sw
tri 38624 25688 38916 25980 ne
rect 38916 25970 42596 25980
tri 42596 25970 42878 26252 sw
tri 42878 25970 43160 26252 ne
rect 43160 26089 46988 26252
tri 46988 26089 47285 26386 sw
tri 47285 26089 47582 26386 ne
rect 47582 26311 49051 26386
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47582 26089 49340 26311
rect 43160 25970 47285 26089
rect 38916 25688 42878 25970
tri 42878 25688 43160 25970 sw
tri 43160 25688 43442 25970 ne
rect 43442 25891 47285 25970
tri 47285 25891 47483 26089 sw
tri 47582 25891 47780 26089 ne
rect 47780 26022 49340 26089
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47780 25891 49629 26022
rect 43442 25688 47483 25891
tri 34380 21444 38624 25688 ne
tri 38624 25396 38916 25688 sw
tri 38916 25396 39208 25688 ne
rect 39208 25406 43160 25688
tri 43160 25406 43442 25688 sw
tri 43442 25406 43724 25688 ne
rect 43724 25594 47483 25688
tri 47483 25594 47780 25891 sw
tri 47780 25594 48077 25891 ne
rect 48077 25778 49629 25891
tri 49629 25778 49873 26022 sw
tri 49918 25778 50162 26022 ne
rect 50162 25778 71000 26022
rect 48077 25594 49873 25778
rect 43724 25406 47780 25594
rect 39208 25396 43442 25406
rect 38624 25104 38916 25396
tri 38916 25104 39208 25396 sw
tri 39208 25104 39500 25396 ne
rect 39500 25208 43442 25396
tri 43442 25208 43640 25406 sw
tri 43724 25208 43922 25406 ne
rect 43922 25297 47780 25406
tri 47780 25297 48077 25594 sw
tri 48077 25297 48374 25594 ne
rect 48374 25489 49873 25594
tri 49873 25489 50162 25778 sw
tri 50162 25489 50451 25778 ne
rect 50451 25489 71000 25778
rect 48374 25297 50162 25489
rect 43922 25208 48077 25297
rect 39500 25104 43640 25208
rect 38624 24812 39208 25104
tri 39208 24812 39500 25104 sw
tri 39500 24812 39792 25104 ne
rect 39792 24926 43640 25104
tri 43640 24926 43922 25208 sw
tri 43922 24926 44204 25208 ne
rect 44204 25000 48077 25208
tri 48077 25000 48374 25297 sw
tri 48374 25000 48671 25297 ne
rect 48671 25200 50162 25297
tri 50162 25200 50451 25489 sw
tri 50451 25200 50740 25489 ne
rect 50740 25200 71000 25489
rect 48671 25000 50451 25200
tri 50451 25000 50651 25200 sw
rect 44204 24926 48374 25000
rect 39792 24812 43922 24926
rect 38624 24520 39500 24812
tri 39500 24520 39792 24812 sw
tri 39792 24520 40084 24812 ne
rect 40084 24644 43922 24812
tri 43922 24644 44204 24926 sw
tri 44204 24644 44486 24926 ne
rect 44486 24703 48374 24926
tri 48374 24703 48671 25000 sw
tri 48671 24703 48968 25000 ne
rect 48968 24906 71000 25000
rect 48968 24703 70613 24906
rect 44486 24644 48671 24703
rect 40084 24520 44204 24644
rect 38624 24228 39792 24520
tri 39792 24228 40084 24520 sw
tri 40084 24228 40376 24520 ne
rect 40376 24362 44204 24520
tri 44204 24362 44486 24644 sw
tri 44486 24362 44768 24644 ne
rect 44768 24406 48671 24644
tri 48671 24406 48968 24703 sw
tri 48968 24406 49265 24703 ne
rect 49265 24406 70613 24703
rect 44768 24362 48968 24406
rect 40376 24228 44486 24362
rect 38624 23948 40084 24228
tri 40084 23948 40364 24228 sw
tri 40376 23948 40656 24228 ne
rect 40656 24080 44486 24228
tri 44486 24080 44768 24362 sw
tri 44768 24080 45050 24362 ne
rect 45050 24194 48968 24362
tri 48968 24194 49180 24406 sw
tri 49265 24194 49477 24406 ne
rect 49477 24194 70613 24406
rect 45050 24080 49180 24194
rect 40656 23948 44768 24080
rect 38624 23656 40364 23948
tri 40364 23656 40656 23948 sw
tri 40656 23656 40948 23948 ne
rect 40948 23798 44768 23948
tri 44768 23798 45050 24080 sw
tri 45050 23798 45332 24080 ne
rect 45332 23897 49180 24080
tri 49180 23897 49477 24194 sw
tri 49477 23897 49774 24194 ne
rect 49774 23897 70613 24194
rect 45332 23798 49477 23897
rect 40948 23656 45050 23798
rect 38624 23364 40656 23656
tri 40656 23364 40948 23656 sw
tri 40948 23364 41240 23656 ne
rect 41240 23516 45050 23656
tri 45050 23516 45332 23798 sw
tri 45332 23516 45614 23798 ne
rect 45614 23600 49477 23798
tri 49477 23600 49774 23897 sw
tri 49774 23600 50071 23897 ne
rect 50071 23706 70613 23897
rect 70669 23706 71000 24906
rect 50071 23600 71000 23706
rect 45614 23516 49774 23600
rect 41240 23364 45332 23516
rect 38624 23072 40948 23364
tri 40948 23072 41240 23364 sw
tri 41240 23072 41532 23364 ne
rect 41532 23234 45332 23364
tri 45332 23234 45614 23516 sw
tri 45614 23234 45896 23516 ne
rect 45896 23400 49774 23516
tri 49774 23400 49974 23600 sw
rect 45896 23234 71000 23400
rect 41532 23072 45614 23234
rect 38624 22780 41240 23072
tri 41240 22780 41532 23072 sw
tri 41532 22780 41824 23072 ne
rect 41824 22952 45614 23072
tri 45614 22952 45896 23234 sw
tri 45896 22952 46178 23234 ne
rect 46178 22952 71000 23234
rect 41824 22854 45896 22952
tri 45896 22854 45994 22952 sw
tri 46178 22854 46276 22952 ne
rect 46276 22854 71000 22952
rect 41824 22780 45994 22854
rect 38624 22488 41532 22780
tri 41532 22488 41824 22780 sw
tri 41824 22488 42116 22780 ne
rect 42116 22572 45994 22780
tri 45994 22572 46276 22854 sw
tri 46276 22572 46558 22854 ne
rect 46558 22572 71000 22854
rect 42116 22488 46276 22572
rect 38624 22196 41824 22488
tri 41824 22196 42116 22488 sw
tri 42116 22196 42408 22488 ne
rect 42408 22290 46276 22488
tri 46276 22290 46558 22572 sw
tri 46558 22290 46840 22572 ne
rect 46840 22290 71000 22572
rect 42408 22196 46558 22290
rect 38624 22028 42116 22196
tri 42116 22028 42284 22196 sw
tri 42408 22028 42576 22196 ne
rect 42576 22028 46558 22196
rect 38624 21736 42284 22028
tri 42284 21736 42576 22028 sw
tri 42576 21736 42868 22028 ne
rect 42868 22008 46558 22028
tri 46558 22008 46840 22290 sw
tri 46840 22008 47122 22290 ne
rect 47122 22008 71000 22290
rect 42868 21736 46840 22008
rect 38624 21444 42576 21736
tri 42576 21444 42868 21736 sw
tri 42868 21444 43160 21736 ne
rect 43160 21726 46840 21736
tri 46840 21726 47122 22008 sw
tri 47122 21726 47404 22008 ne
rect 47404 21726 71000 22008
rect 43160 21444 47122 21726
tri 47122 21444 47404 21726 sw
tri 47404 21444 47686 21726 ne
rect 47686 21444 71000 21726
tri 38624 17200 42868 21444 ne
tri 42868 21152 43160 21444 sw
tri 43160 21152 43452 21444 ne
rect 43452 21162 47404 21444
tri 47404 21162 47686 21444 sw
tri 47686 21162 47968 21444 ne
rect 47968 21162 71000 21444
rect 43452 21152 47686 21162
rect 42868 20860 43160 21152
tri 43160 20860 43452 21152 sw
tri 43452 20860 43744 21152 ne
rect 43744 20964 47686 21152
tri 47686 20964 47884 21162 sw
tri 47968 20964 48166 21162 ne
rect 48166 20964 71000 21162
rect 43744 20860 47884 20964
rect 42868 20568 43452 20860
tri 43452 20568 43744 20860 sw
tri 43744 20568 44036 20860 ne
rect 44036 20682 47884 20860
tri 47884 20682 48166 20964 sw
tri 48166 20682 48448 20964 ne
rect 48448 20682 71000 20964
rect 44036 20568 48166 20682
rect 42868 20276 43744 20568
tri 43744 20276 44036 20568 sw
tri 44036 20276 44328 20568 ne
rect 44328 20400 48166 20568
tri 48166 20400 48448 20682 sw
tri 48448 20400 48730 20682 ne
rect 48730 20400 71000 20682
rect 44328 20276 48448 20400
rect 42868 19984 44036 20276
tri 44036 19984 44328 20276 sw
tri 44328 19984 44620 20276 ne
rect 44620 20200 48448 20276
tri 48448 20200 48648 20400 sw
rect 44620 19984 71000 20200
rect 42868 19704 44328 19984
tri 44328 19704 44608 19984 sw
tri 44620 19704 44900 19984 ne
rect 44900 19704 71000 19984
rect 42868 19412 44608 19704
tri 44608 19412 44900 19704 sw
tri 44900 19412 45192 19704 ne
rect 45192 19412 71000 19704
rect 42868 19120 44900 19412
tri 44900 19120 45192 19412 sw
tri 45192 19120 45484 19412 ne
rect 45484 19120 71000 19412
rect 42868 18828 45192 19120
tri 45192 18828 45484 19120 sw
tri 45484 18828 45776 19120 ne
rect 45776 18828 71000 19120
rect 42868 18536 45484 18828
tri 45484 18536 45776 18828 sw
tri 45776 18536 46068 18828 ne
rect 46068 18536 71000 18828
rect 42868 18244 45776 18536
tri 45776 18244 46068 18536 sw
tri 46068 18244 46360 18536 ne
rect 46360 18244 71000 18536
rect 42868 17952 46068 18244
tri 46068 17952 46360 18244 sw
tri 46360 17952 46652 18244 ne
rect 46652 17952 71000 18244
rect 42868 17784 46360 17952
tri 46360 17784 46528 17952 sw
tri 46652 17784 46820 17952 ne
rect 46820 17784 71000 17952
rect 42868 17492 46528 17784
tri 46528 17492 46820 17784 sw
tri 46820 17492 47112 17784 ne
rect 47112 17492 71000 17784
rect 42868 17200 46820 17492
tri 46820 17200 47112 17492 sw
tri 47112 17200 47404 17492 ne
rect 47404 17200 71000 17492
tri 42868 14000 46068 17200 ne
rect 46068 17000 47112 17200
tri 47112 17000 47312 17200 sw
rect 46068 14000 71000 17000
<< labels >>
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 1 nsew
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 1 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 2 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 2 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 3 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 4 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 4 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 4 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 4 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 4 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 4 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 4 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 4 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 4 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 4 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 4 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string GDS_END 29533672
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 28534372
<< end >>
