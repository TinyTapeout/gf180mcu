magic
tech gf180mcuD
magscale 1 10
timestamp 1764353313
<< nwell >>
rect 361 13779 14639 69307
<< obsm1 >>
rect -32 13108 15032 69957
<< metal2 >>
rect 672 65709 748 70000
rect 1193 66084 1269 70000
rect 1422 65374 1498 70000
rect 1564 65256 1640 70001
rect 2066 66020 2142 70000
rect 2277 66984 2353 70000
rect 13734 53268 13810 70000
rect 13880 53414 13956 70000
rect 14026 56689 14102 70000
rect 14172 63980 14248 70000
<< obsm2 >>
rect 0 65649 612 69675
rect 808 66024 1133 69675
rect 1329 66024 1362 69675
rect 808 65649 1362 66024
rect 0 65314 1362 65649
rect 0 65196 1504 65314
rect 1700 65960 2006 69675
rect 2202 66924 2217 69675
rect 2413 66924 13674 69675
rect 2202 65960 13674 66924
rect 1700 65196 13674 65960
rect 0 53208 13674 65196
rect 14308 63920 15000 69675
rect 14162 56629 15000 63920
rect 14016 53354 15000 56629
rect 13870 53208 15000 53354
rect 0 0 15000 53208
<< obsm3 >>
rect 0 0 15000 69678
<< obsm4 >>
rect 0 0 15000 69678
<< metal5 >>
rect 0 68400 1000 69678
rect 0 66800 1000 68200
rect 0 65200 1000 66600
rect 0 63600 1000 65000
rect 0 62000 1000 63400
rect 0 60400 1000 61800
rect 0 58800 1000 60200
rect 0 57200 1000 58600
rect 0 55600 1000 57000
rect 0 54000 1000 55400
rect 0 52400 1000 53800
rect 0 50800 1000 52200
rect 0 49200 1000 50600
rect 0 46000 1000 49000
rect 0 42800 1000 45800
rect 0 41200 1000 42600
rect 0 39600 1000 41000
rect 0 36400 1000 39400
rect 0 33200 1000 36200
rect 0 30000 1000 33000
rect 0 26800 1000 29800
rect 0 25200 1000 26600
rect 0 23600 1000 25000
rect 0 20400 1000 23400
rect 0 17200 1000 20200
rect 0 14000 1000 17000
rect 14000 68400 15000 69678
rect 14000 66800 15000 68200
rect 14000 65200 15000 66600
rect 14000 63600 15000 65000
rect 14000 62000 15000 63400
rect 14000 60400 15000 61800
rect 14000 58800 15000 60200
rect 14000 57200 15000 58600
rect 14000 55600 15000 57000
rect 14000 54000 15000 55400
rect 14000 52400 15000 53800
rect 14000 50800 15000 52200
rect 14000 49200 15000 50600
rect 14000 46000 15000 49000
rect 14000 42800 15000 45800
rect 14000 41200 15000 42600
rect 14000 39600 15000 41000
rect 14000 36400 15000 39400
rect 14000 33200 15000 36200
rect 14000 30000 15000 33000
rect 14000 26800 15000 29800
rect 14000 25200 15000 26600
rect 14000 23600 15000 25000
rect 14000 20400 15000 23400
rect 14000 17200 15000 20200
rect 14000 14000 15000 17000
rect 1500 400 13500 12400
<< obsm5 >>
rect 1120 13880 13880 69678
rect 700 12520 14300 13880
rect 700 280 1380 12520
rect 13620 280 14300 12520
rect 700 0 14300 280
<< labels >>
rlabel metal2 s 13880 53414 13956 70000 6 A
port 1 nsew signal input
rlabel metal2 s 672 65709 748 70000 6 CS
port 2 nsew signal input
rlabel metal5 s 0 36400 1000 39400 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 42800 1000 45800 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 66800 1000 68200 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 58800 1000 60200 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 55600 1000 57000 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 54000 1000 55400 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 52400 1000 53800 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 41200 1000 42600 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 23600 1000 25000 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 26800 1000 29800 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 30000 1000 33000 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 33200 1000 36200 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 36400 15000 39400 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 42800 15000 45800 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 66800 15000 68200 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 58800 15000 60200 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 55600 15000 57000 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 54000 15000 55400 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 52400 15000 53800 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 41200 15000 42600 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 23600 15000 25000 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 26800 15000 29800 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 30000 15000 33000 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 14000 33200 15000 36200 6 DVDD
port 3 nsew power bidirectional
rlabel metal5 s 0 17200 1000 20200 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 14000 1000 17000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 46000 1000 49000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 39600 1000 41000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 20400 1000 23400 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 25200 1000 26600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 57200 1000 58600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 60400 1000 61800 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 65200 1000 66600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 68400 1000 69678 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 17200 15000 20200 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 14000 15000 17000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 46000 15000 49000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 39600 15000 41000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 20400 15000 23400 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 25200 15000 26600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 57200 15000 58600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 60400 15000 61800 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 65200 15000 66600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal5 s 14000 68400 15000 69678 6 DVSS
port 4 nsew ground bidirectional
rlabel metal2 s 2277 66984 2353 70000 6 IE
port 5 nsew signal input
rlabel metal2 s 14026 56689 14102 70000 6 OE
port 6 nsew signal input
rlabel metal5 s 1500 400 13500 12400 6 PAD
port 7 nsew signal bidirectional
rlabel metal2 s 2066 66020 2142 70000 6 PD
port 8 nsew signal input
rlabel metal2 s 1422 65374 1498 70000 6 PDRV0
port 9 nsew signal input
rlabel metal2 s 1564 65256 1640 70001 6 PDRV1
port 10 nsew signal input
rlabel metal2 s 1193 66084 1269 70000 6 PU
port 11 nsew signal input
rlabel metal2 s 13734 53268 13810 70000 6 SL
port 12 nsew signal input
rlabel metal5 s 0 50800 1000 52200 6 VDD
port 13 nsew power bidirectional
rlabel metal5 s 0 62000 1000 63400 6 VDD
port 13 nsew power bidirectional
rlabel metal5 s 14000 50800 15000 52200 6 VDD
port 13 nsew power bidirectional
rlabel metal5 s 14000 62000 15000 63400 6 VDD
port 13 nsew power bidirectional
rlabel metal5 s 0 63600 1000 65000 6 VSS
port 14 nsew ground bidirectional
rlabel metal5 s 0 49200 1000 50600 6 VSS
port 14 nsew ground bidirectional
rlabel metal5 s 14000 63600 15000 65000 6 VSS
port 14 nsew ground bidirectional
rlabel metal5 s 14000 49200 15000 50600 6 VSS
port 14 nsew ground bidirectional
rlabel metal2 s 14172 63980 14248 70000 6 Y
port 15 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string LEFclass PAD INOUT
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 13940822
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_ocd_io/gds/gf180mcu_ocd_io.gds
string GDS_START 13928198
<< end >>
